module tt_um_Samcooper01 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \curr_seg[0] ;
 wire \curr_seg[1] ;
 wire \curr_seg[2] ;
 wire \curr_seg[3] ;
 wire \feistel_out_q[0] ;
 wire \feistel_out_q[1] ;
 wire \feistel_out_q[2] ;
 wire \feistel_out_q[3] ;
 wire \feistel_out_q[4] ;
 wire \feistel_out_q[5] ;
 wire \feistel_out_q[6] ;
 wire \feistel_out_q[7] ;
 wire \key_bytes[0][4] ;
 wire \key_bytes[0][5] ;
 wire \key_bytes[0][6] ;
 wire \key_bytes[0][7] ;
 wire \key_bytes[10][4] ;
 wire \key_bytes[10][5] ;
 wire \key_bytes[10][6] ;
 wire \key_bytes[10][7] ;
 wire \key_bytes[11][4] ;
 wire \key_bytes[11][5] ;
 wire \key_bytes[11][6] ;
 wire \key_bytes[11][7] ;
 wire \key_bytes[12][4] ;
 wire \key_bytes[12][5] ;
 wire \key_bytes[12][6] ;
 wire \key_bytes[12][7] ;
 wire \key_bytes[13][4] ;
 wire \key_bytes[13][5] ;
 wire \key_bytes[13][6] ;
 wire \key_bytes[13][7] ;
 wire \key_bytes[14][4] ;
 wire \key_bytes[14][5] ;
 wire \key_bytes[14][6] ;
 wire \key_bytes[14][7] ;
 wire \key_bytes[15][4] ;
 wire \key_bytes[15][5] ;
 wire \key_bytes[15][6] ;
 wire \key_bytes[15][7] ;
 wire \key_bytes[1][4] ;
 wire \key_bytes[1][5] ;
 wire \key_bytes[1][6] ;
 wire \key_bytes[1][7] ;
 wire \key_bytes[2][4] ;
 wire \key_bytes[2][5] ;
 wire \key_bytes[2][6] ;
 wire \key_bytes[2][7] ;
 wire \key_bytes[3][4] ;
 wire \key_bytes[3][5] ;
 wire \key_bytes[3][6] ;
 wire \key_bytes[3][7] ;
 wire \key_bytes[4][4] ;
 wire \key_bytes[4][5] ;
 wire \key_bytes[4][6] ;
 wire \key_bytes[4][7] ;
 wire \key_bytes[5][4] ;
 wire \key_bytes[5][5] ;
 wire \key_bytes[5][6] ;
 wire \key_bytes[5][7] ;
 wire \key_bytes[6][4] ;
 wire \key_bytes[6][5] ;
 wire \key_bytes[6][6] ;
 wire \key_bytes[6][7] ;
 wire \key_bytes[7][4] ;
 wire \key_bytes[7][5] ;
 wire \key_bytes[7][6] ;
 wire \key_bytes[7][7] ;
 wire \key_bytes[8][4] ;
 wire \key_bytes[8][5] ;
 wire \key_bytes[8][6] ;
 wire \key_bytes[8][7] ;
 wire \key_bytes[9][4] ;
 wire \key_bytes[9][5] ;
 wire \key_bytes[9][6] ;
 wire \key_bytes[9][7] ;
 wire mode_dec;
 wire out_valid;
 wire prev_streaming;
 wire \start_seg[0] ;
 wire \start_seg[1] ;
 wire \start_seg[2] ;
 wire \start_seg[3] ;
 wire \sys_next_state[0] ;
 wire \sys_next_state[1] ;
 wire \sys_state[0] ;
 wire \sys_state[1] ;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;

 sky130_fd_sc_hd__inv_2 _0478_ (.A(net3),
    .Y(_0085_));
 sky130_fd_sc_hd__inv_2 _0479_ (.A(\start_seg[2] ),
    .Y(_0086_));
 sky130_fd_sc_hd__inv_2 _0480_ (.A(net31),
    .Y(_0087_));
 sky130_fd_sc_hd__and2_1 _0481_ (.A(\sys_state[0] ),
    .B(net22),
    .X(_0477_));
 sky130_fd_sc_hd__nand2b_1 _0482_ (.A_N(net22),
    .B(\sys_state[0] ),
    .Y(_0088_));
 sky130_fd_sc_hd__nor2_1 _0483_ (.A(net134),
    .B(_0088_),
    .Y(_0000_));
 sky130_fd_sc_hd__nand2_2 _0484_ (.A(\counter[1] ),
    .B(_0000_),
    .Y(_0089_));
 sky130_fd_sc_hd__or3b_4 _0485_ (.A(\counter[1] ),
    .B(_0088_),
    .C_N(\counter[0] ),
    .X(_0090_));
 sky130_fd_sc_hd__nand2_1 _0486_ (.A(_0089_),
    .B(_0090_),
    .Y(_0001_));
 sky130_fd_sc_hd__and3_1 _0487_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .C(\counter[2] ),
    .X(_0091_));
 sky130_fd_sc_hd__a21oi_1 _0488_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .B1(\counter[2] ),
    .Y(_0092_));
 sky130_fd_sc_hd__nor3_1 _0489_ (.A(_0088_),
    .B(_0091_),
    .C(_0092_),
    .Y(_0002_));
 sky130_fd_sc_hd__nand2_1 _0490_ (.A(\counter[2] ),
    .B(\counter[3] ),
    .Y(_0093_));
 sky130_fd_sc_hd__a21oi_1 _0491_ (.A1(\counter[3] ),
    .A2(_0091_),
    .B1(_0088_),
    .Y(_0094_));
 sky130_fd_sc_hd__o21a_1 _0492_ (.A1(\counter[3] ),
    .A2(_0091_),
    .B1(_0094_),
    .X(_0003_));
 sky130_fd_sc_hd__nor4b_1 _0493_ (.A(net29),
    .B(net27),
    .C(net23),
    .D_N(net25),
    .Y(_0095_));
 sky130_fd_sc_hd__and4bb_1 _0494_ (.A_N(net27),
    .B_N(net26),
    .C(net24),
    .D(net29),
    .X(_0096_));
 sky130_fd_sc_hd__a22o_1 _0495_ (.A1(\key_bytes[4][5] ),
    .A2(net20),
    .B1(_0096_),
    .B2(\key_bytes[9][5] ),
    .X(_0097_));
 sky130_fd_sc_hd__and4_1 _0496_ (.A(net30),
    .B(net27),
    .C(net25),
    .D(net23),
    .X(_0098_));
 sky130_fd_sc_hd__and4b_2 _0497_ (.A_N(net23),
    .B(net25),
    .C(net28),
    .D(net30),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_1 _0498_ (.A1(\key_bytes[15][5] ),
    .A2(_0098_),
    .B1(_0099_),
    .B2(\key_bytes[7][5] ),
    .X(_0100_));
 sky130_fd_sc_hd__or4_4 _0499_ (.A(\curr_seg[0] ),
    .B(net28),
    .C(net26),
    .D(net24),
    .X(_0101_));
 sky130_fd_sc_hd__and4b_1 _0500_ (.A_N(net29),
    .B(net28),
    .C(net26),
    .D(net24),
    .X(_0102_));
 sky130_fd_sc_hd__a21bo_1 _0501_ (.A1(\key_bytes[14][5] ),
    .A2(_0102_),
    .B1_N(_0101_),
    .X(_0103_));
 sky130_fd_sc_hd__and4bb_1 _0502_ (.A_N(net30),
    .B_N(net23),
    .C(net25),
    .D(net27),
    .X(_0104_));
 sky130_fd_sc_hd__and4b_1 _0503_ (.A_N(net27),
    .B(net25),
    .C(net23),
    .D(net30),
    .X(_0105_));
 sky130_fd_sc_hd__a22o_1 _0504_ (.A1(\key_bytes[6][5] ),
    .A2(_0104_),
    .B1(_0105_),
    .B2(\key_bytes[13][5] ),
    .X(_0106_));
 sky130_fd_sc_hd__or4_1 _0505_ (.A(_0097_),
    .B(_0100_),
    .C(_0103_),
    .D(_0106_),
    .X(_0107_));
 sky130_fd_sc_hd__and4bb_1 _0506_ (.A_N(net26),
    .B_N(net24),
    .C(net29),
    .D(net28),
    .X(_0108_));
 sky130_fd_sc_hd__and4b_1 _0507_ (.A_N(net26),
    .B(net24),
    .C(net29),
    .D(net28),
    .X(_0109_));
 sky130_fd_sc_hd__a22o_1 _0508_ (.A1(\key_bytes[3][5] ),
    .A2(_0108_),
    .B1(_0109_),
    .B2(\key_bytes[11][5] ),
    .X(_0110_));
 sky130_fd_sc_hd__and4bb_2 _0509_ (.A_N(net30),
    .B_N(\curr_seg[1] ),
    .C(net26),
    .D(net24),
    .X(_0111_));
 sky130_fd_sc_hd__and4bb_1 _0510_ (.A_N(net27),
    .B_N(net23),
    .C(net25),
    .D(net29),
    .X(_0112_));
 sky130_fd_sc_hd__a22o_1 _0511_ (.A1(\key_bytes[12][5] ),
    .A2(_0111_),
    .B1(_0112_),
    .B2(\key_bytes[5][5] ),
    .X(_0113_));
 sky130_fd_sc_hd__nor4b_1 _0512_ (.A(net27),
    .B(net25),
    .C(net23),
    .D_N(net29),
    .Y(_0114_));
 sky130_fd_sc_hd__nor4b_1 _0513_ (.A(net29),
    .B(net27),
    .C(net25),
    .D_N(net23),
    .Y(_0115_));
 sky130_fd_sc_hd__a22o_1 _0514_ (.A1(\key_bytes[1][5] ),
    .A2(net19),
    .B1(net18),
    .B2(\key_bytes[8][5] ),
    .X(_0116_));
 sky130_fd_sc_hd__nor4b_1 _0515_ (.A(net29),
    .B(net26),
    .C(net24),
    .D_N(net28),
    .Y(_0117_));
 sky130_fd_sc_hd__and4bb_1 _0516_ (.A_N(net29),
    .B_N(net25),
    .C(net23),
    .D(net27),
    .X(_0118_));
 sky130_fd_sc_hd__a22o_1 _0517_ (.A1(\key_bytes[2][5] ),
    .A2(net17),
    .B1(_0118_),
    .B2(\key_bytes[10][5] ),
    .X(_0119_));
 sky130_fd_sc_hd__or4_1 _0518_ (.A(_0110_),
    .B(_0113_),
    .C(_0116_),
    .D(_0119_),
    .X(_0120_));
 sky130_fd_sc_hd__or2_1 _0519_ (.A(\key_bytes[0][5] ),
    .B(_0101_),
    .X(_0121_));
 sky130_fd_sc_hd__and3_2 _0520_ (.A(\sys_state[0] ),
    .B(net22),
    .C(net47),
    .X(_0122_));
 sky130_fd_sc_hd__o211a_1 _0521_ (.A1(_0107_),
    .A2(_0120_),
    .B1(_0121_),
    .C1(_0122_),
    .X(_0123_));
 sky130_fd_sc_hd__xnor2_4 _0522_ (.A(\start_seg[1] ),
    .B(_0123_),
    .Y(_0124_));
 sky130_fd_sc_hd__inv_2 _0523_ (.A(_0124_),
    .Y(_0125_));
 sky130_fd_sc_hd__a22o_1 _0524_ (.A1(\key_bytes[9][4] ),
    .A2(_0096_),
    .B1(_0112_),
    .B2(\key_bytes[5][4] ),
    .X(_0126_));
 sky130_fd_sc_hd__a22o_1 _0525_ (.A1(\key_bytes[15][4] ),
    .A2(_0098_),
    .B1(net18),
    .B2(\key_bytes[8][4] ),
    .X(_0127_));
 sky130_fd_sc_hd__a21bo_1 _0526_ (.A1(\key_bytes[13][4] ),
    .A2(_0105_),
    .B1_N(_0101_),
    .X(_0128_));
 sky130_fd_sc_hd__a22o_1 _0527_ (.A1(\key_bytes[7][4] ),
    .A2(_0099_),
    .B1(_0111_),
    .B2(\key_bytes[12][4] ),
    .X(_0129_));
 sky130_fd_sc_hd__or4_1 _0528_ (.A(_0126_),
    .B(_0127_),
    .C(_0128_),
    .D(_0129_),
    .X(_0130_));
 sky130_fd_sc_hd__a22o_1 _0529_ (.A1(\key_bytes[14][4] ),
    .A2(_0102_),
    .B1(_0117_),
    .B2(\key_bytes[2][4] ),
    .X(_0131_));
 sky130_fd_sc_hd__a22o_1 _0530_ (.A1(\key_bytes[6][4] ),
    .A2(_0104_),
    .B1(_0118_),
    .B2(\key_bytes[10][4] ),
    .X(_0132_));
 sky130_fd_sc_hd__a22o_1 _0531_ (.A1(\key_bytes[4][4] ),
    .A2(net20),
    .B1(_0114_),
    .B2(\key_bytes[1][4] ),
    .X(_0133_));
 sky130_fd_sc_hd__a22o_1 _0532_ (.A1(\key_bytes[3][4] ),
    .A2(_0108_),
    .B1(_0109_),
    .B2(\key_bytes[11][4] ),
    .X(_0134_));
 sky130_fd_sc_hd__or4_1 _0533_ (.A(_0131_),
    .B(_0132_),
    .C(_0133_),
    .D(_0134_),
    .X(_0135_));
 sky130_fd_sc_hd__or2_1 _0534_ (.A(\key_bytes[0][4] ),
    .B(_0101_),
    .X(_0136_));
 sky130_fd_sc_hd__o211a_1 _0535_ (.A1(_0130_),
    .A2(_0135_),
    .B1(_0136_),
    .C1(_0122_),
    .X(_0137_));
 sky130_fd_sc_hd__xor2_2 _0536_ (.A(\start_seg[0] ),
    .B(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__xnor2_1 _0537_ (.A(\start_seg[0] ),
    .B(_0137_),
    .Y(_0139_));
 sky130_fd_sc_hd__a22o_1 _0538_ (.A1(\key_bytes[9][6] ),
    .A2(_0096_),
    .B1(net17),
    .B2(\key_bytes[2][6] ),
    .X(_0140_));
 sky130_fd_sc_hd__a22o_1 _0539_ (.A1(\key_bytes[14][6] ),
    .A2(_0102_),
    .B1(_0109_),
    .B2(\key_bytes[11][6] ),
    .X(_0141_));
 sky130_fd_sc_hd__a21bo_1 _0540_ (.A1(\key_bytes[12][6] ),
    .A2(_0111_),
    .B1_N(_0101_),
    .X(_0142_));
 sky130_fd_sc_hd__a22o_1 _0541_ (.A1(\key_bytes[4][6] ),
    .A2(net20),
    .B1(_0108_),
    .B2(\key_bytes[3][6] ),
    .X(_0143_));
 sky130_fd_sc_hd__or4_1 _0542_ (.A(_0140_),
    .B(_0141_),
    .C(_0142_),
    .D(_0143_),
    .X(_0144_));
 sky130_fd_sc_hd__a22o_1 _0543_ (.A1(\key_bytes[8][6] ),
    .A2(net18),
    .B1(_0118_),
    .B2(\key_bytes[10][6] ),
    .X(_0145_));
 sky130_fd_sc_hd__a221o_1 _0544_ (.A1(\key_bytes[15][6] ),
    .A2(_0098_),
    .B1(_0105_),
    .B2(\key_bytes[13][6] ),
    .C1(_0145_),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _0545_ (.A1(\key_bytes[6][6] ),
    .A2(_0104_),
    .B1(_0112_),
    .B2(\key_bytes[5][6] ),
    .X(_0147_));
 sky130_fd_sc_hd__a221o_1 _0546_ (.A1(\key_bytes[7][6] ),
    .A2(_0099_),
    .B1(net19),
    .B2(\key_bytes[1][6] ),
    .C1(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__nor3_2 _0547_ (.A(_0144_),
    .B(_0146_),
    .C(_0148_),
    .Y(_0149_));
 sky130_fd_sc_hd__o21ai_2 _0548_ (.A1(\key_bytes[0][6] ),
    .A2(_0101_),
    .B1(_0122_),
    .Y(_0150_));
 sky130_fd_sc_hd__or3_2 _0549_ (.A(_0086_),
    .B(_0149_),
    .C(_0150_),
    .X(_0151_));
 sky130_fd_sc_hd__o21ai_4 _0550_ (.A1(_0149_),
    .A2(_0150_),
    .B1(_0086_),
    .Y(_0152_));
 sky130_fd_sc_hd__nand2_4 _0551_ (.A(_0151_),
    .B(_0152_),
    .Y(_0153_));
 sky130_fd_sc_hd__nand2_1 _0552_ (.A(\start_seg[0] ),
    .B(\start_seg[1] ),
    .Y(_0154_));
 sky130_fd_sc_hd__nand3_1 _0553_ (.A(_0151_),
    .B(_0152_),
    .C(_0154_),
    .Y(_0155_));
 sky130_fd_sc_hd__a21o_1 _0554_ (.A1(_0151_),
    .A2(_0152_),
    .B1(_0154_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_2 _0555_ (.A(_0155_),
    .B(_0156_),
    .X(_0157_));
 sky130_fd_sc_hd__nand3_2 _0556_ (.A(net4),
    .B(_0151_),
    .C(_0152_),
    .Y(_0158_));
 sky130_fd_sc_hd__a21o_1 _0557_ (.A1(_0151_),
    .A2(_0152_),
    .B1(net4),
    .X(_0159_));
 sky130_fd_sc_hd__nand2_1 _0558_ (.A(_0085_),
    .B(_0124_),
    .Y(_0160_));
 sky130_fd_sc_hd__a2bb2o_1 _0559_ (.A1_N(_0085_),
    .A2_N(_0124_),
    .B1(_0138_),
    .B2(net42),
    .X(_0161_));
 sky130_fd_sc_hd__nand4_2 _0560_ (.A(_0158_),
    .B(_0159_),
    .C(_0160_),
    .D(_0161_),
    .Y(_0162_));
 sky130_fd_sc_hd__a22o_1 _0561_ (.A1(_0158_),
    .A2(_0159_),
    .B1(_0160_),
    .B2(_0161_),
    .X(_0163_));
 sky130_fd_sc_hd__xnor2_1 _0562_ (.A(net3),
    .B(net36),
    .Y(_0164_));
 sky130_fd_sc_hd__nand3_1 _0563_ (.A(_0162_),
    .B(_0163_),
    .C(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__a21o_1 _0564_ (.A1(_0162_),
    .A2(_0163_),
    .B1(_0164_),
    .X(_0166_));
 sky130_fd_sc_hd__nand2_1 _0565_ (.A(_0165_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__a21o_1 _0566_ (.A1(_0165_),
    .A2(_0166_),
    .B1(_0157_),
    .X(_0168_));
 sky130_fd_sc_hd__nand3_1 _0567_ (.A(_0157_),
    .B(_0165_),
    .C(_0166_),
    .Y(_0169_));
 sky130_fd_sc_hd__xnor2_1 _0568_ (.A(\start_seg[0] ),
    .B(_0124_),
    .Y(_0170_));
 sky130_fd_sc_hd__inv_2 _0569_ (.A(net13),
    .Y(_0171_));
 sky130_fd_sc_hd__xnor2_1 _0570_ (.A(net3),
    .B(_0124_),
    .Y(_0172_));
 sky130_fd_sc_hd__or3b_1 _0571_ (.A(net38),
    .B(net16),
    .C_N(net42),
    .X(_0173_));
 sky130_fd_sc_hd__a21bo_1 _0572_ (.A1(net42),
    .A2(net15),
    .B1_N(net38),
    .X(_0174_));
 sky130_fd_sc_hd__nand2_1 _0573_ (.A(_0173_),
    .B(_0174_),
    .Y(_0175_));
 sky130_fd_sc_hd__a21oi_1 _0574_ (.A1(_0173_),
    .A2(_0174_),
    .B1(_0172_),
    .Y(_0176_));
 sky130_fd_sc_hd__and3_1 _0575_ (.A(_0172_),
    .B(_0173_),
    .C(_0174_),
    .X(_0177_));
 sky130_fd_sc_hd__nor2_1 _0576_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__nand2_1 _0577_ (.A(net40),
    .B(net16),
    .Y(_0179_));
 sky130_fd_sc_hd__xnor2_1 _0578_ (.A(net40),
    .B(net16),
    .Y(_0180_));
 sky130_fd_sc_hd__xor2_1 _0579_ (.A(net42),
    .B(net5),
    .X(_0181_));
 sky130_fd_sc_hd__xnor2_1 _0580_ (.A(_0180_),
    .B(_0181_),
    .Y(_0182_));
 sky130_fd_sc_hd__o31a_1 _0581_ (.A1(net13),
    .A2(_0176_),
    .A3(_0177_),
    .B1(_0182_),
    .X(_0183_));
 sky130_fd_sc_hd__a2bb2o_1 _0582_ (.A1_N(_0171_),
    .A2_N(_0178_),
    .B1(_0183_),
    .B2(net15),
    .X(_0184_));
 sky130_fd_sc_hd__nand3_1 _0583_ (.A(_0168_),
    .B(_0169_),
    .C(_0184_),
    .Y(_0185_));
 sky130_fd_sc_hd__nand2_2 _0584_ (.A(_0168_),
    .B(_0185_),
    .Y(_0186_));
 sky130_fd_sc_hd__nand2_2 _0585_ (.A(\start_seg[2] ),
    .B(\start_seg[1] ),
    .Y(_0187_));
 sky130_fd_sc_hd__a22o_1 _0586_ (.A1(\key_bytes[5][7] ),
    .A2(_0112_),
    .B1(net19),
    .B2(\key_bytes[1][7] ),
    .X(_0188_));
 sky130_fd_sc_hd__a22o_1 _0587_ (.A1(\key_bytes[3][7] ),
    .A2(_0108_),
    .B1(_0109_),
    .B2(\key_bytes[11][7] ),
    .X(_0189_));
 sky130_fd_sc_hd__a221o_1 _0588_ (.A1(\key_bytes[14][7] ),
    .A2(_0102_),
    .B1(_0117_),
    .B2(\key_bytes[2][7] ),
    .C1(_0189_),
    .X(_0190_));
 sky130_fd_sc_hd__a211o_1 _0589_ (.A1(\key_bytes[15][7] ),
    .A2(_0098_),
    .B1(_0188_),
    .C1(_0190_),
    .X(_0191_));
 sky130_fd_sc_hd__a22o_1 _0590_ (.A1(\key_bytes[9][7] ),
    .A2(_0096_),
    .B1(_0099_),
    .B2(\key_bytes[7][7] ),
    .X(_0192_));
 sky130_fd_sc_hd__a221o_1 _0591_ (.A1(\key_bytes[4][7] ),
    .A2(_0095_),
    .B1(_0115_),
    .B2(\key_bytes[8][7] ),
    .C1(_0192_),
    .X(_0193_));
 sky130_fd_sc_hd__a22o_1 _0592_ (.A1(\key_bytes[12][7] ),
    .A2(_0111_),
    .B1(_0118_),
    .B2(\key_bytes[10][7] ),
    .X(_0194_));
 sky130_fd_sc_hd__a21bo_1 _0593_ (.A1(\key_bytes[6][7] ),
    .A2(_0104_),
    .B1_N(_0101_),
    .X(_0195_));
 sky130_fd_sc_hd__a2111o_1 _0594_ (.A1(\key_bytes[13][7] ),
    .A2(_0105_),
    .B1(_0193_),
    .C1(_0194_),
    .D1(_0195_),
    .X(_0196_));
 sky130_fd_sc_hd__o221ai_4 _0595_ (.A1(\key_bytes[0][7] ),
    .A2(_0101_),
    .B1(_0191_),
    .B2(_0196_),
    .C1(_0122_),
    .Y(_0197_));
 sky130_fd_sc_hd__xor2_4 _0596_ (.A(\start_seg[3] ),
    .B(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__xnor2_4 _0597_ (.A(_0187_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__mux2_2 _0598_ (.A0(net12),
    .A1(_0199_),
    .S(\start_seg[0] ),
    .X(_0200_));
 sky130_fd_sc_hd__nand2_2 _0599_ (.A(_0158_),
    .B(_0162_),
    .Y(_0201_));
 sky130_fd_sc_hd__nor2_1 _0600_ (.A(net4),
    .B(net5),
    .Y(_0202_));
 sky130_fd_sc_hd__and2_1 _0601_ (.A(net4),
    .B(net5),
    .X(_0203_));
 sky130_fd_sc_hd__nor2_1 _0602_ (.A(_0202_),
    .B(_0203_),
    .Y(_0204_));
 sky130_fd_sc_hd__xnor2_1 _0603_ (.A(net34),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__xnor2_2 _0604_ (.A(_0198_),
    .B(_0205_),
    .Y(_0206_));
 sky130_fd_sc_hd__xnor2_4 _0605_ (.A(_0201_),
    .B(_0206_),
    .Y(_0207_));
 sky130_fd_sc_hd__xnor2_1 _0606_ (.A(_0200_),
    .B(_0207_),
    .Y(_0208_));
 sky130_fd_sc_hd__xnor2_1 _0607_ (.A(net5),
    .B(_0167_),
    .Y(_0209_));
 sky130_fd_sc_hd__xnor2_2 _0608_ (.A(_0208_),
    .B(_0209_),
    .Y(_0210_));
 sky130_fd_sc_hd__xor2_4 _0609_ (.A(_0186_),
    .B(_0210_),
    .X(_0211_));
 sky130_fd_sc_hd__xor2_1 _0610_ (.A(net42),
    .B(_0207_),
    .X(_0212_));
 sky130_fd_sc_hd__xnor2_2 _0611_ (.A(_0211_),
    .B(_0212_),
    .Y(_0213_));
 sky130_fd_sc_hd__nand2_2 _0612_ (.A(net16),
    .B(_0213_),
    .Y(_0214_));
 sky130_fd_sc_hd__nand2_2 _0613_ (.A(_0138_),
    .B(_0182_),
    .Y(_0215_));
 sky130_fd_sc_hd__xnor2_2 _0614_ (.A(\start_seg[0] ),
    .B(_0175_),
    .Y(_0216_));
 sky130_fd_sc_hd__xnor2_4 _0615_ (.A(_0215_),
    .B(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__xnor2_2 _0616_ (.A(net5),
    .B(net41),
    .Y(_0218_));
 sky130_fd_sc_hd__xnor2_4 _0617_ (.A(_0207_),
    .B(_0218_),
    .Y(_0219_));
 sky130_fd_sc_hd__or2_2 _0618_ (.A(_0138_),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__xnor2_1 _0619_ (.A(_0124_),
    .B(_0217_),
    .Y(_0221_));
 sky130_fd_sc_hd__xnor2_2 _0620_ (.A(_0178_),
    .B(_0221_),
    .Y(_0222_));
 sky130_fd_sc_hd__xnor2_4 _0621_ (.A(_0220_),
    .B(_0222_),
    .Y(_0223_));
 sky130_fd_sc_hd__xnor2_1 _0622_ (.A(net13),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__xnor2_2 _0623_ (.A(_0217_),
    .B(_0224_),
    .Y(_0225_));
 sky130_fd_sc_hd__xor2_4 _0624_ (.A(_0214_),
    .B(_0225_),
    .X(_0226_));
 sky130_fd_sc_hd__a21o_1 _0625_ (.A1(_0168_),
    .A2(_0169_),
    .B1(_0184_),
    .X(_0227_));
 sky130_fd_sc_hd__xnor2_1 _0626_ (.A(net4),
    .B(_0178_),
    .Y(_0228_));
 sky130_fd_sc_hd__nand3_1 _0627_ (.A(_0185_),
    .B(_0227_),
    .C(_0228_),
    .Y(_0229_));
 sky130_fd_sc_hd__a21o_1 _0628_ (.A1(_0185_),
    .A2(_0227_),
    .B1(_0228_),
    .X(_0230_));
 sky130_fd_sc_hd__nand2_1 _0629_ (.A(_0229_),
    .B(_0230_),
    .Y(_0231_));
 sky130_fd_sc_hd__xnor2_2 _0630_ (.A(\start_seg[1] ),
    .B(_0153_),
    .Y(_0232_));
 sky130_fd_sc_hd__nand3_1 _0631_ (.A(_0229_),
    .B(_0230_),
    .C(_0232_),
    .Y(_0233_));
 sky130_fd_sc_hd__a211o_1 _0632_ (.A1(_0125_),
    .A2(_0217_),
    .B1(_0219_),
    .C1(net15),
    .X(_0234_));
 sky130_fd_sc_hd__o21ai_1 _0633_ (.A1(_0125_),
    .A2(_0217_),
    .B1(_0234_),
    .Y(_0235_));
 sky130_fd_sc_hd__a21o_1 _0634_ (.A1(_0229_),
    .A2(_0230_),
    .B1(_0232_),
    .X(_0236_));
 sky130_fd_sc_hd__nand3_1 _0635_ (.A(_0233_),
    .B(_0235_),
    .C(_0236_),
    .Y(_0237_));
 sky130_fd_sc_hd__a21boi_1 _0636_ (.A1(_0235_),
    .A2(_0236_),
    .B1_N(_0233_),
    .Y(_0238_));
 sky130_fd_sc_hd__xnor2_1 _0637_ (.A(_0207_),
    .B(_0231_),
    .Y(_0239_));
 sky130_fd_sc_hd__xor2_1 _0638_ (.A(_0199_),
    .B(_0211_),
    .X(_0240_));
 sky130_fd_sc_hd__xnor2_1 _0639_ (.A(_0238_),
    .B(_0240_),
    .Y(_0241_));
 sky130_fd_sc_hd__xnor2_1 _0640_ (.A(_0239_),
    .B(_0241_),
    .Y(_0242_));
 sky130_fd_sc_hd__xnor2_1 _0641_ (.A(_0219_),
    .B(_0242_),
    .Y(_0243_));
 sky130_fd_sc_hd__or2_1 _0642_ (.A(_0138_),
    .B(_0213_),
    .X(_0244_));
 sky130_fd_sc_hd__and2_1 _0643_ (.A(_0214_),
    .B(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__xnor2_1 _0644_ (.A(_0243_),
    .B(_0245_),
    .Y(_0246_));
 sky130_fd_sc_hd__a21oi_1 _0645_ (.A1(_0124_),
    .A2(_0226_),
    .B1(net15),
    .Y(_0247_));
 sky130_fd_sc_hd__o2bb2a_1 _0646_ (.A1_N(_0247_),
    .A2_N(_0246_),
    .B1(_0226_),
    .B2(_0124_),
    .X(_0248_));
 sky130_fd_sc_hd__nor2_2 _0647_ (.A(\start_seg[0] ),
    .B(\start_seg[1] ),
    .Y(_0249_));
 sky130_fd_sc_hd__xor2_2 _0648_ (.A(_0153_),
    .B(_0249_),
    .X(_0250_));
 sky130_fd_sc_hd__xnor2_1 _0649_ (.A(_0153_),
    .B(_0249_),
    .Y(_0251_));
 sky130_fd_sc_hd__a21o_1 _0650_ (.A1(_0233_),
    .A2(_0236_),
    .B1(_0235_),
    .X(_0252_));
 sky130_fd_sc_hd__xnor2_1 _0651_ (.A(_0167_),
    .B(_0217_),
    .Y(_0253_));
 sky130_fd_sc_hd__nand3_1 _0652_ (.A(_0237_),
    .B(_0252_),
    .C(_0253_),
    .Y(_0254_));
 sky130_fd_sc_hd__a21o_1 _0653_ (.A1(_0237_),
    .A2(_0252_),
    .B1(_0253_),
    .X(_0255_));
 sky130_fd_sc_hd__nand2_1 _0654_ (.A(_0254_),
    .B(_0255_),
    .Y(_0256_));
 sky130_fd_sc_hd__nand3_1 _0655_ (.A(_0250_),
    .B(_0254_),
    .C(_0255_),
    .Y(_0257_));
 sky130_fd_sc_hd__a21o_1 _0656_ (.A1(_0254_),
    .A2(_0255_),
    .B1(_0250_),
    .X(_0258_));
 sky130_fd_sc_hd__o211a_1 _0657_ (.A1(_0171_),
    .A2(_0223_),
    .B1(_0213_),
    .C1(net15),
    .X(_0259_));
 sky130_fd_sc_hd__a21o_1 _0658_ (.A1(_0171_),
    .A2(_0223_),
    .B1(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__nand3_1 _0659_ (.A(_0257_),
    .B(_0258_),
    .C(_0260_),
    .Y(_0261_));
 sky130_fd_sc_hd__a21o_1 _0660_ (.A1(_0257_),
    .A2(_0258_),
    .B1(_0260_),
    .X(_0262_));
 sky130_fd_sc_hd__xor2_1 _0661_ (.A(_0223_),
    .B(_0231_),
    .X(_0263_));
 sky130_fd_sc_hd__a21o_1 _0662_ (.A1(_0261_),
    .A2(_0262_),
    .B1(_0263_),
    .X(_0264_));
 sky130_fd_sc_hd__nand3_1 _0663_ (.A(_0261_),
    .B(_0262_),
    .C(_0263_),
    .Y(_0265_));
 sky130_fd_sc_hd__nand2_1 _0664_ (.A(_0264_),
    .B(_0265_),
    .Y(_0266_));
 sky130_fd_sc_hd__a21o_1 _0665_ (.A1(_0264_),
    .A2(_0265_),
    .B1(_0153_),
    .X(_0267_));
 sky130_fd_sc_hd__nand3_1 _0666_ (.A(_0153_),
    .B(_0264_),
    .C(_0265_),
    .Y(_0268_));
 sky130_fd_sc_hd__mux2_1 _0667_ (.A0(_0268_),
    .A1(_0267_),
    .S(_0248_),
    .X(_0269_));
 sky130_fd_sc_hd__nand2_2 _0668_ (.A(_0257_),
    .B(_0261_),
    .Y(_0270_));
 sky130_fd_sc_hd__nor2_2 _0669_ (.A(_0086_),
    .B(_0249_),
    .Y(_0271_));
 sky130_fd_sc_hd__xnor2_4 _0670_ (.A(net12),
    .B(_0271_),
    .Y(_0272_));
 sky130_fd_sc_hd__xnor2_1 _0671_ (.A(_0211_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__xnor2_2 _0672_ (.A(_0256_),
    .B(_0273_),
    .Y(_0274_));
 sky130_fd_sc_hd__xnor2_4 _0673_ (.A(_0270_),
    .B(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__xnor2_2 _0674_ (.A(\start_seg[2] ),
    .B(_0198_),
    .Y(_0276_));
 sky130_fd_sc_hd__xnor2_1 _0675_ (.A(_0242_),
    .B(_0275_),
    .Y(_0277_));
 sky130_fd_sc_hd__xor2_1 _0676_ (.A(_0275_),
    .B(_0276_),
    .X(_0278_));
 sky130_fd_sc_hd__xnor2_2 _0677_ (.A(_0269_),
    .B(_0278_),
    .Y(_0279_));
 sky130_fd_sc_hd__xnor2_1 _0678_ (.A(_0213_),
    .B(_0277_),
    .Y(_0280_));
 sky130_fd_sc_hd__nor2_1 _0679_ (.A(_0279_),
    .B(_0280_),
    .Y(_0281_));
 sky130_fd_sc_hd__a21o_1 _0680_ (.A1(_0279_),
    .A2(_0280_),
    .B1(net31),
    .X(_0282_));
 sky130_fd_sc_hd__and3_1 _0681_ (.A(net35),
    .B(_0155_),
    .C(_0156_),
    .X(_0283_));
 sky130_fd_sc_hd__a21o_1 _0682_ (.A1(_0155_),
    .A2(_0156_),
    .B1(net35),
    .X(_0284_));
 sky130_fd_sc_hd__and2b_1 _0683_ (.A_N(_0283_),
    .B(_0284_),
    .X(_0285_));
 sky130_fd_sc_hd__or2_1 _0684_ (.A(net37),
    .B(net13),
    .X(_0286_));
 sky130_fd_sc_hd__nand2_1 _0685_ (.A(net37),
    .B(net13),
    .Y(_0287_));
 sky130_fd_sc_hd__a22o_1 _0686_ (.A1(net40),
    .A2(net14),
    .B1(net13),
    .B2(net37),
    .X(_0288_));
 sky130_fd_sc_hd__nand2_1 _0687_ (.A(_0286_),
    .B(_0288_),
    .Y(_0289_));
 sky130_fd_sc_hd__xnor2_1 _0688_ (.A(_0285_),
    .B(_0289_),
    .Y(_0290_));
 sky130_fd_sc_hd__xor2_1 _0689_ (.A(net4),
    .B(net37),
    .X(_0291_));
 sky130_fd_sc_hd__xnor2_1 _0690_ (.A(_0290_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__or2_1 _0691_ (.A(_0153_),
    .B(_0292_),
    .X(_0293_));
 sky130_fd_sc_hd__nand2_1 _0692_ (.A(_0153_),
    .B(_0292_),
    .Y(_0294_));
 sky130_fd_sc_hd__nand2_1 _0693_ (.A(_0293_),
    .B(_0294_),
    .Y(_0295_));
 sky130_fd_sc_hd__xnor2_2 _0694_ (.A(_0085_),
    .B(_0179_),
    .Y(_0296_));
 sky130_fd_sc_hd__a21oi_1 _0695_ (.A1(_0286_),
    .A2(_0287_),
    .B1(_0296_),
    .Y(_0297_));
 sky130_fd_sc_hd__and3_1 _0696_ (.A(_0286_),
    .B(_0287_),
    .C(_0296_),
    .X(_0298_));
 sky130_fd_sc_hd__or2_2 _0697_ (.A(_0297_),
    .B(_0298_),
    .X(_0299_));
 sky130_fd_sc_hd__xnor2_2 _0698_ (.A(net42),
    .B(net33),
    .Y(_0300_));
 sky130_fd_sc_hd__xnor2_1 _0699_ (.A(_0180_),
    .B(_0300_),
    .Y(_0301_));
 sky130_fd_sc_hd__xnor2_1 _0700_ (.A(net35),
    .B(_0299_),
    .Y(_0302_));
 sky130_fd_sc_hd__o211a_1 _0701_ (.A1(_0125_),
    .A2(_0299_),
    .B1(_0301_),
    .C1(net16),
    .X(_0303_));
 sky130_fd_sc_hd__a21o_1 _0702_ (.A1(_0125_),
    .A2(_0299_),
    .B1(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__xnor2_1 _0703_ (.A(_0302_),
    .B(_0304_),
    .Y(_0305_));
 sky130_fd_sc_hd__xnor2_2 _0704_ (.A(_0295_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__xnor2_1 _0705_ (.A(_0250_),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__nand2_2 _0706_ (.A(net14),
    .B(_0301_),
    .Y(_0308_));
 sky130_fd_sc_hd__xnor2_2 _0707_ (.A(\start_seg[0] ),
    .B(_0296_),
    .Y(_0309_));
 sky130_fd_sc_hd__xnor2_4 _0708_ (.A(_0308_),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__a31o_1 _0709_ (.A1(_0284_),
    .A2(_0286_),
    .A3(_0288_),
    .B1(_0283_),
    .X(_0311_));
 sky130_fd_sc_hd__and2_1 _0710_ (.A(_0086_),
    .B(_0154_),
    .X(_0312_));
 sky130_fd_sc_hd__xnor2_2 _0711_ (.A(net12),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__xor2_1 _0712_ (.A(net33),
    .B(net36),
    .X(_0314_));
 sky130_fd_sc_hd__xnor2_1 _0713_ (.A(net5),
    .B(_0314_),
    .Y(_0315_));
 sky130_fd_sc_hd__xnor2_2 _0714_ (.A(_0313_),
    .B(_0315_),
    .Y(_0316_));
 sky130_fd_sc_hd__xnor2_2 _0715_ (.A(_0311_),
    .B(_0316_),
    .Y(_0317_));
 sky130_fd_sc_hd__xnor2_1 _0716_ (.A(_0300_),
    .B(_0317_),
    .Y(_0318_));
 sky130_fd_sc_hd__o21bai_1 _0717_ (.A1(_0171_),
    .A2(_0310_),
    .B1_N(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__o2bb2a_1 _0718_ (.A1_N(_0171_),
    .A2_N(_0310_),
    .B1(_0319_),
    .B2(net16),
    .X(_0320_));
 sky130_fd_sc_hd__xnor2_1 _0719_ (.A(_0307_),
    .B(_0320_),
    .Y(_0321_));
 sky130_fd_sc_hd__xnor2_1 _0720_ (.A(_0292_),
    .B(_0310_),
    .Y(_0322_));
 sky130_fd_sc_hd__xnor2_2 _0721_ (.A(_0321_),
    .B(_0322_),
    .Y(_0323_));
 sky130_fd_sc_hd__nor2_2 _0722_ (.A(net14),
    .B(_0318_),
    .Y(_0324_));
 sky130_fd_sc_hd__xnor2_1 _0723_ (.A(_0171_),
    .B(_0310_),
    .Y(_0325_));
 sky130_fd_sc_hd__xnor2_2 _0724_ (.A(_0299_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__xnor2_4 _0725_ (.A(_0324_),
    .B(_0326_),
    .Y(_0327_));
 sky130_fd_sc_hd__xor2_2 _0726_ (.A(net33),
    .B(_0276_),
    .X(_0328_));
 sky130_fd_sc_hd__mux2_1 _0727_ (.A0(_0293_),
    .A1(_0294_),
    .S(_0304_),
    .X(_0329_));
 sky130_fd_sc_hd__xnor2_2 _0728_ (.A(_0328_),
    .B(_0329_),
    .Y(_0330_));
 sky130_fd_sc_hd__xor2_2 _0729_ (.A(net40),
    .B(_0330_),
    .X(_0331_));
 sky130_fd_sc_hd__a21o_1 _0730_ (.A1(_0125_),
    .A2(_0327_),
    .B1(net14),
    .X(_0332_));
 sky130_fd_sc_hd__o22ai_1 _0731_ (.A1(_0125_),
    .A2(_0327_),
    .B1(_0331_),
    .B2(_0332_),
    .Y(_0333_));
 sky130_fd_sc_hd__nor2_1 _0732_ (.A(_0232_),
    .B(_0333_),
    .Y(_0334_));
 sky130_fd_sc_hd__and2_1 _0733_ (.A(_0232_),
    .B(_0333_),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_1 _0734_ (.A0(_0334_),
    .A1(_0335_),
    .S(_0323_),
    .X(_0336_));
 sky130_fd_sc_hd__xnor2_2 _0735_ (.A(_0199_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__xor2_1 _0736_ (.A(_0300_),
    .B(_0330_),
    .X(_0338_));
 sky130_fd_sc_hd__xnor2_2 _0737_ (.A(_0337_),
    .B(_0338_),
    .Y(_0339_));
 sky130_fd_sc_hd__o221a_1 _0738_ (.A1(_0281_),
    .A2(_0282_),
    .B1(_0339_),
    .B2(_0087_),
    .C1(net21),
    .X(_0004_));
 sky130_fd_sc_hd__xnor2_2 _0739_ (.A(_0219_),
    .B(_0275_),
    .Y(_0340_));
 sky130_fd_sc_hd__inv_2 _0740_ (.A(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__nand2_2 _0741_ (.A(net15),
    .B(_0246_),
    .Y(_0342_));
 sky130_fd_sc_hd__xnor2_1 _0742_ (.A(_0124_),
    .B(_0226_),
    .Y(_0343_));
 sky130_fd_sc_hd__xnor2_2 _0743_ (.A(_0223_),
    .B(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__xnor2_4 _0744_ (.A(_0342_),
    .B(_0344_),
    .Y(_0345_));
 sky130_fd_sc_hd__xnor2_1 _0745_ (.A(_0171_),
    .B(_0345_),
    .Y(_0346_));
 sky130_fd_sc_hd__xnor2_1 _0746_ (.A(_0226_),
    .B(_0346_),
    .Y(_0347_));
 sky130_fd_sc_hd__or3_1 _0747_ (.A(net14),
    .B(_0340_),
    .C(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__o21ai_1 _0748_ (.A1(net14),
    .A2(_0340_),
    .B1(_0347_),
    .Y(_0349_));
 sky130_fd_sc_hd__xor2_1 _0749_ (.A(_0272_),
    .B(_0330_),
    .X(_0350_));
 sky130_fd_sc_hd__mux2_1 _0750_ (.A0(_0251_),
    .A1(_0306_),
    .S(_0320_),
    .X(_0351_));
 sky130_fd_sc_hd__o21ba_1 _0751_ (.A1(_0251_),
    .A2(_0306_),
    .B1_N(_0351_),
    .X(_0352_));
 sky130_fd_sc_hd__xnor2_1 _0752_ (.A(_0350_),
    .B(_0352_),
    .Y(_0353_));
 sky130_fd_sc_hd__and2_1 _0753_ (.A(net14),
    .B(_0318_),
    .X(_0354_));
 sky130_fd_sc_hd__nor2_1 _0754_ (.A(_0324_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__xnor2_1 _0755_ (.A(_0331_),
    .B(_0355_),
    .Y(_0356_));
 sky130_fd_sc_hd__xor2_1 _0756_ (.A(_0353_),
    .B(_0356_),
    .X(_0357_));
 sky130_fd_sc_hd__nor2_1 _0757_ (.A(net14),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__nor2_2 _0758_ (.A(net16),
    .B(_0331_),
    .Y(_0359_));
 sky130_fd_sc_hd__xnor2_1 _0759_ (.A(_0124_),
    .B(_0327_),
    .Y(_0360_));
 sky130_fd_sc_hd__xnor2_2 _0760_ (.A(_0310_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__xnor2_4 _0761_ (.A(_0359_),
    .B(_0361_),
    .Y(_0362_));
 sky130_fd_sc_hd__nand2_1 _0762_ (.A(net13),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__nor2_1 _0763_ (.A(net13),
    .B(_0362_),
    .Y(_0364_));
 sky130_fd_sc_hd__xnor2_1 _0764_ (.A(net13),
    .B(_0362_),
    .Y(_0365_));
 sky130_fd_sc_hd__xnor2_1 _0765_ (.A(_0327_),
    .B(_0365_),
    .Y(_0366_));
 sky130_fd_sc_hd__xnor2_2 _0766_ (.A(_0358_),
    .B(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__o21ai_1 _0767_ (.A1(_0087_),
    .A2(_0367_),
    .B1(net21),
    .Y(_0368_));
 sky130_fd_sc_hd__a31oi_1 _0768_ (.A1(_0087_),
    .A2(_0348_),
    .A3(_0349_),
    .B1(_0368_),
    .Y(_0005_));
 sky130_fd_sc_hd__xor2_1 _0769_ (.A(_0226_),
    .B(_0256_),
    .X(_0369_));
 sky130_fd_sc_hd__inv_2 _0770_ (.A(_0369_),
    .Y(_0370_));
 sky130_fd_sc_hd__and3_1 _0771_ (.A(_0248_),
    .B(_0267_),
    .C(_0268_),
    .X(_0371_));
 sky130_fd_sc_hd__a21oi_1 _0772_ (.A1(_0267_),
    .A2(_0268_),
    .B1(_0248_),
    .Y(_0372_));
 sky130_fd_sc_hd__or3_1 _0773_ (.A(_0370_),
    .B(_0371_),
    .C(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__o21ai_1 _0774_ (.A1(_0371_),
    .A2(_0372_),
    .B1(_0370_),
    .Y(_0374_));
 sky130_fd_sc_hd__and2_1 _0775_ (.A(_0373_),
    .B(_0374_),
    .X(_0375_));
 sky130_fd_sc_hd__and3_1 _0776_ (.A(_0157_),
    .B(_0373_),
    .C(_0374_),
    .X(_0376_));
 sky130_fd_sc_hd__a21o_1 _0777_ (.A1(_0373_),
    .A2(_0374_),
    .B1(_0157_),
    .X(_0377_));
 sky130_fd_sc_hd__nand2b_1 _0778_ (.A_N(_0376_),
    .B(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__a2bb2o_1 _0779_ (.A1_N(net16),
    .A2_N(_0340_),
    .B1(_0345_),
    .B2(net13),
    .X(_0379_));
 sky130_fd_sc_hd__o21a_1 _0780_ (.A1(_0170_),
    .A2(_0345_),
    .B1(_0379_),
    .X(_0380_));
 sky130_fd_sc_hd__xnor2_1 _0781_ (.A(_0378_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__xnor2_1 _0782_ (.A(_0266_),
    .B(_0345_),
    .Y(_0382_));
 sky130_fd_sc_hd__xnor2_1 _0783_ (.A(_0381_),
    .B(_0382_),
    .Y(_0383_));
 sky130_fd_sc_hd__or2_1 _0784_ (.A(_0334_),
    .B(_0335_),
    .X(_0384_));
 sky130_fd_sc_hd__xnor2_1 _0785_ (.A(_0306_),
    .B(_0327_),
    .Y(_0385_));
 sky130_fd_sc_hd__xnor2_1 _0786_ (.A(_0323_),
    .B(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__xnor2_2 _0787_ (.A(_0384_),
    .B(_0386_),
    .Y(_0387_));
 sky130_fd_sc_hd__nor2_1 _0788_ (.A(_0157_),
    .B(_0387_),
    .Y(_0388_));
 sky130_fd_sc_hd__and2_1 _0789_ (.A(_0157_),
    .B(_0387_),
    .X(_0389_));
 sky130_fd_sc_hd__or2_1 _0790_ (.A(_0388_),
    .B(_0389_),
    .X(_0390_));
 sky130_fd_sc_hd__o31a_1 _0791_ (.A1(net16),
    .A2(_0357_),
    .A3(_0364_),
    .B1(_0363_),
    .X(_0391_));
 sky130_fd_sc_hd__xnor2_1 _0792_ (.A(_0390_),
    .B(_0391_),
    .Y(_0392_));
 sky130_fd_sc_hd__xor2_1 _0793_ (.A(_0323_),
    .B(_0362_),
    .X(_0393_));
 sky130_fd_sc_hd__xnor2_1 _0794_ (.A(_0392_),
    .B(_0393_),
    .Y(_0394_));
 sky130_fd_sc_hd__nand2_1 _0795_ (.A(net31),
    .B(_0394_),
    .Y(_0395_));
 sky130_fd_sc_hd__o211a_1 _0796_ (.A1(net31),
    .A2(_0383_),
    .B1(_0395_),
    .C1(net21),
    .X(_0006_));
 sky130_fd_sc_hd__a21oi_1 _0797_ (.A1(_0377_),
    .A2(_0380_),
    .B1(_0376_),
    .Y(_0396_));
 sky130_fd_sc_hd__xnor2_1 _0798_ (.A(_0277_),
    .B(_0396_),
    .Y(_0397_));
 sky130_fd_sc_hd__xor2_1 _0799_ (.A(_0279_),
    .B(_0313_),
    .X(_0398_));
 sky130_fd_sc_hd__nor2_1 _0800_ (.A(_0375_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__a31o_1 _0801_ (.A1(_0373_),
    .A2(_0374_),
    .A3(_0398_),
    .B1(_0399_),
    .X(_0400_));
 sky130_fd_sc_hd__nor2_1 _0802_ (.A(_0397_),
    .B(_0400_),
    .Y(_0401_));
 sky130_fd_sc_hd__a21o_1 _0803_ (.A1(_0397_),
    .A2(_0400_),
    .B1(mode_dec),
    .X(_0402_));
 sky130_fd_sc_hd__o21bai_2 _0804_ (.A1(_0390_),
    .A2(_0391_),
    .B1_N(_0388_),
    .Y(_0403_));
 sky130_fd_sc_hd__xnor2_1 _0805_ (.A(_0272_),
    .B(_0317_),
    .Y(_0404_));
 sky130_fd_sc_hd__xnor2_1 _0806_ (.A(_0352_),
    .B(_0404_),
    .Y(_0405_));
 sky130_fd_sc_hd__xnor2_1 _0807_ (.A(_0337_),
    .B(_0405_),
    .Y(_0406_));
 sky130_fd_sc_hd__xor2_1 _0808_ (.A(_0200_),
    .B(_0353_),
    .X(_0407_));
 sky130_fd_sc_hd__xnor2_1 _0809_ (.A(_0387_),
    .B(_0407_),
    .Y(_0408_));
 sky130_fd_sc_hd__xnor2_1 _0810_ (.A(_0406_),
    .B(_0408_),
    .Y(_0409_));
 sky130_fd_sc_hd__xnor2_2 _0811_ (.A(_0403_),
    .B(_0409_),
    .Y(_0410_));
 sky130_fd_sc_hd__nand2_1 _0812_ (.A(net31),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__o211a_1 _0813_ (.A1(_0401_),
    .A2(_0402_),
    .B1(_0411_),
    .C1(_0477_),
    .X(_0007_));
 sky130_fd_sc_hd__and2_1 _0814_ (.A(net14),
    .B(_0357_),
    .X(_0412_));
 sky130_fd_sc_hd__or2_1 _0815_ (.A(_0358_),
    .B(_0412_),
    .X(_0413_));
 sky130_fd_sc_hd__xnor2_1 _0816_ (.A(_0339_),
    .B(_0413_),
    .Y(_0414_));
 sky130_fd_sc_hd__nor2_1 _0817_ (.A(_0410_),
    .B(_0414_),
    .Y(_0415_));
 sky130_fd_sc_hd__a21o_1 _0818_ (.A1(_0410_),
    .A2(_0414_),
    .B1(_0087_),
    .X(_0416_));
 sky130_fd_sc_hd__o221a_1 _0819_ (.A1(mode_dec),
    .A2(_0341_),
    .B1(_0415_),
    .B2(_0416_),
    .C1(net21),
    .X(_0008_));
 sky130_fd_sc_hd__or2_1 _0820_ (.A(_0125_),
    .B(_0367_),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _0821_ (.A(_0125_),
    .B(_0367_),
    .Y(_0418_));
 sky130_fd_sc_hd__and2_1 _0822_ (.A(_0417_),
    .B(_0418_),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_1 _0823_ (.A(net14),
    .B(_0339_),
    .Y(_0420_));
 sky130_fd_sc_hd__xor2_1 _0824_ (.A(_0362_),
    .B(_0420_),
    .X(_0421_));
 sky130_fd_sc_hd__and2_1 _0825_ (.A(_0419_),
    .B(_0421_),
    .X(_0422_));
 sky130_fd_sc_hd__o21ai_1 _0826_ (.A1(_0419_),
    .A2(_0421_),
    .B1(net31),
    .Y(_0423_));
 sky130_fd_sc_hd__o221a_1 _0827_ (.A1(net31),
    .A2(_0345_),
    .B1(_0422_),
    .B2(_0423_),
    .C1(net21),
    .X(_0009_));
 sky130_fd_sc_hd__xor2_1 _0828_ (.A(_0367_),
    .B(_0387_),
    .X(_0424_));
 sky130_fd_sc_hd__o211ai_1 _0829_ (.A1(_0125_),
    .A2(_0367_),
    .B1(_0339_),
    .C1(net16),
    .Y(_0425_));
 sky130_fd_sc_hd__and3_1 _0830_ (.A(_0153_),
    .B(_0418_),
    .C(_0425_),
    .X(_0426_));
 sky130_fd_sc_hd__a21oi_1 _0831_ (.A1(_0418_),
    .A2(_0425_),
    .B1(_0153_),
    .Y(_0427_));
 sky130_fd_sc_hd__nor2_1 _0832_ (.A(_0426_),
    .B(_0427_),
    .Y(_0428_));
 sky130_fd_sc_hd__xnor2_1 _0833_ (.A(_0394_),
    .B(_0428_),
    .Y(_0429_));
 sky130_fd_sc_hd__nor2_1 _0834_ (.A(_0424_),
    .B(_0429_),
    .Y(_0430_));
 sky130_fd_sc_hd__a21o_1 _0835_ (.A1(_0424_),
    .A2(_0429_),
    .B1(_0087_),
    .X(_0431_));
 sky130_fd_sc_hd__o221a_1 _0836_ (.A1(net31),
    .A2(_0375_),
    .B1(_0430_),
    .B2(_0431_),
    .C1(net21),
    .X(_0010_));
 sky130_fd_sc_hd__xnor2_1 _0837_ (.A(net12),
    .B(_0408_),
    .Y(_0432_));
 sky130_fd_sc_hd__xnor2_1 _0838_ (.A(_0403_),
    .B(_0432_),
    .Y(_0433_));
 sky130_fd_sc_hd__mux2_1 _0839_ (.A0(_0426_),
    .A1(_0427_),
    .S(_0394_),
    .X(_0434_));
 sky130_fd_sc_hd__nor2_1 _0840_ (.A(_0433_),
    .B(_0434_),
    .Y(_0435_));
 sky130_fd_sc_hd__a21o_1 _0841_ (.A1(_0433_),
    .A2(_0434_),
    .B1(_0087_),
    .X(_0436_));
 sky130_fd_sc_hd__o221a_1 _0842_ (.A1(net31),
    .A2(_0279_),
    .B1(_0435_),
    .B2(_0436_),
    .C1(net21),
    .X(_0011_));
 sky130_fd_sc_hd__or4_1 _0843_ (.A(net41),
    .B(net34),
    .C(net36),
    .D(net38),
    .X(_0437_));
 sky130_fd_sc_hd__nor2_1 _0844_ (.A(\sys_state[0] ),
    .B(net22),
    .Y(_0438_));
 sky130_fd_sc_hd__nand2_1 _0845_ (.A(_0202_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__and2_1 _0846_ (.A(net42),
    .B(net3),
    .X(_0440_));
 sky130_fd_sc_hd__nor2_1 _0847_ (.A(net42),
    .B(net3),
    .Y(_0441_));
 sky130_fd_sc_hd__and2b_1 _0848_ (.A_N(net11),
    .B(net21),
    .X(_0442_));
 sky130_fd_sc_hd__or4_1 _0849_ (.A(_0437_),
    .B(_0439_),
    .C(_0440_),
    .D(_0441_),
    .X(_0443_));
 sky130_fd_sc_hd__or3b_1 _0850_ (.A(_0094_),
    .B(_0442_),
    .C_N(_0443_),
    .X(\sys_next_state[0] ));
 sky130_fd_sc_hd__mux2_1 _0851_ (.A0(_0202_),
    .A1(_0203_),
    .S(net2),
    .X(_0444_));
 sky130_fd_sc_hd__nor2_1 _0852_ (.A(_0085_),
    .B(_0437_),
    .Y(_0445_));
 sky130_fd_sc_hd__a31o_1 _0853_ (.A1(_0438_),
    .A2(_0444_),
    .A3(_0445_),
    .B1(_0442_),
    .X(\sys_next_state[1] ));
 sky130_fd_sc_hd__and2_2 _0854_ (.A(out_valid),
    .B(\feistel_out_q[0] ),
    .X(uo_out[0]));
 sky130_fd_sc_hd__and2_2 _0855_ (.A(out_valid),
    .B(\feistel_out_q[1] ),
    .X(uo_out[1]));
 sky130_fd_sc_hd__and2_2 _0856_ (.A(out_valid),
    .B(\feistel_out_q[2] ),
    .X(uo_out[2]));
 sky130_fd_sc_hd__and2_2 _0857_ (.A(out_valid),
    .B(\feistel_out_q[3] ),
    .X(uo_out[3]));
 sky130_fd_sc_hd__and2_2 _0858_ (.A(out_valid),
    .B(\feistel_out_q[4] ),
    .X(uo_out[4]));
 sky130_fd_sc_hd__and2_2 _0859_ (.A(out_valid),
    .B(\feistel_out_q[5] ),
    .X(uo_out[5]));
 sky130_fd_sc_hd__and2_2 _0860_ (.A(out_valid),
    .B(\feistel_out_q[6] ),
    .X(uo_out[6]));
 sky130_fd_sc_hd__and2_2 _0861_ (.A(out_valid),
    .B(\feistel_out_q[7] ),
    .X(uo_out[7]));
 sky130_fd_sc_hd__mux2_1 _0862_ (.A0(net10),
    .A1(net31),
    .S(net21),
    .X(_0012_));
 sky130_fd_sc_hd__nand2_1 _0863_ (.A(net30),
    .B(_0477_),
    .Y(_0446_));
 sky130_fd_sc_hd__and2b_1 _0864_ (.A_N(\sys_state[0] ),
    .B(\sys_state[1] ),
    .X(_0447_));
 sky130_fd_sc_hd__nand2b_2 _0865_ (.A_N(\sys_state[0] ),
    .B(net22),
    .Y(_0448_));
 sky130_fd_sc_hd__o221a_1 _0866_ (.A1(net22),
    .A2(net30),
    .B1(net42),
    .B2(_0448_),
    .C1(_0446_),
    .X(_0013_));
 sky130_fd_sc_hd__xor2_1 _0867_ (.A(net30),
    .B(net28),
    .X(_0449_));
 sky130_fd_sc_hd__and2b_1 _0868_ (.A_N(\sys_state[1] ),
    .B(net28),
    .X(_0450_));
 sky130_fd_sc_hd__a221o_1 _0869_ (.A1(net3),
    .A2(_0447_),
    .B1(_0449_),
    .B2(net21),
    .C1(_0450_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _0870_ (.A(net4),
    .B(_0447_),
    .X(_0451_));
 sky130_fd_sc_hd__a31o_1 _0871_ (.A1(net22),
    .A2(\curr_seg[0] ),
    .A3(net27),
    .B1(net25),
    .X(_0452_));
 sky130_fd_sc_hd__nand4_1 _0872_ (.A(net22),
    .B(net30),
    .C(net28),
    .D(net26),
    .Y(_0453_));
 sky130_fd_sc_hd__a31o_1 _0873_ (.A1(_0448_),
    .A2(_0452_),
    .A3(_0453_),
    .B1(_0451_),
    .X(_0015_));
 sky130_fd_sc_hd__a21o_1 _0874_ (.A1(net23),
    .A2(_0453_),
    .B1(_0099_),
    .X(_0454_));
 sky130_fd_sc_hd__mux2_1 _0875_ (.A0(net24),
    .A1(\sys_state[0] ),
    .S(net22),
    .X(_0455_));
 sky130_fd_sc_hd__a22o_1 _0876_ (.A1(net5),
    .A2(_0447_),
    .B1(_0454_),
    .B2(_0455_),
    .X(_0016_));
 sky130_fd_sc_hd__and4b_2 _0877_ (.A_N(net22),
    .B(\counter[0] ),
    .C(\counter[1] ),
    .D(\sys_state[0] ),
    .X(_0456_));
 sky130_fd_sc_hd__nand2b_2 _0878_ (.A_N(_0093_),
    .B(_0456_),
    .Y(_0457_));
 sky130_fd_sc_hd__mux2_1 _0879_ (.A0(net39),
    .A1(net120),
    .S(_0457_),
    .X(_0017_));
 sky130_fd_sc_hd__mux2_1 _0880_ (.A0(net38),
    .A1(net71),
    .S(_0457_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0881_ (.A0(net36),
    .A1(net133),
    .S(_0457_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0882_ (.A0(net33),
    .A1(\key_bytes[0][7] ),
    .S(_0457_),
    .X(_0020_));
 sky130_fd_sc_hd__nor2_2 _0883_ (.A(_0089_),
    .B(_0093_),
    .Y(_0458_));
 sky130_fd_sc_hd__mux2_1 _0884_ (.A0(net94),
    .A1(net39),
    .S(_0458_),
    .X(_0021_));
 sky130_fd_sc_hd__mux2_1 _0885_ (.A0(net119),
    .A1(net37),
    .S(_0458_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0886_ (.A0(net114),
    .A1(net35),
    .S(_0458_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0887_ (.A0(net128),
    .A1(net32),
    .S(_0458_),
    .X(_0024_));
 sky130_fd_sc_hd__nor2_1 _0888_ (.A(_0090_),
    .B(_0093_),
    .Y(_0459_));
 sky130_fd_sc_hd__mux2_1 _0889_ (.A0(net77),
    .A1(net41),
    .S(_0459_),
    .X(_0025_));
 sky130_fd_sc_hd__mux2_1 _0890_ (.A0(net91),
    .A1(net38),
    .S(_0459_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _0891_ (.A0(net84),
    .A1(net36),
    .S(_0459_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _0892_ (.A0(net80),
    .A1(net34),
    .S(_0459_),
    .X(_0028_));
 sky130_fd_sc_hd__or3_2 _0893_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .C(_0088_),
    .X(_0460_));
 sky130_fd_sc_hd__nor2_1 _0894_ (.A(_0093_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__mux2_1 _0895_ (.A0(net118),
    .A1(net41),
    .S(_0461_),
    .X(_0029_));
 sky130_fd_sc_hd__mux2_1 _0896_ (.A0(net100),
    .A1(net38),
    .S(_0461_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _0897_ (.A0(net109),
    .A1(net36),
    .S(_0461_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _0898_ (.A0(net106),
    .A1(net34),
    .S(_0461_),
    .X(_0032_));
 sky130_fd_sc_hd__nand2b_2 _0899_ (.A_N(\counter[2] ),
    .B(\counter[3] ),
    .Y(_0462_));
 sky130_fd_sc_hd__nand3b_2 _0900_ (.A_N(\counter[2] ),
    .B(\counter[3] ),
    .C(_0456_),
    .Y(_0463_));
 sky130_fd_sc_hd__mux2_1 _0901_ (.A0(net39),
    .A1(net101),
    .S(_0463_),
    .X(_0033_));
 sky130_fd_sc_hd__mux2_1 _0902_ (.A0(net38),
    .A1(net104),
    .S(_0463_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _0903_ (.A0(net36),
    .A1(net116),
    .S(_0463_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _0904_ (.A0(net32),
    .A1(net115),
    .S(_0463_),
    .X(_0036_));
 sky130_fd_sc_hd__nor2_2 _0905_ (.A(_0089_),
    .B(_0462_),
    .Y(_0464_));
 sky130_fd_sc_hd__mux2_1 _0906_ (.A0(net110),
    .A1(net39),
    .S(_0464_),
    .X(_0037_));
 sky130_fd_sc_hd__mux2_1 _0907_ (.A0(net90),
    .A1(net37),
    .S(_0464_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _0908_ (.A0(net121),
    .A1(net35),
    .S(_0464_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _0909_ (.A0(net87),
    .A1(net32),
    .S(_0464_),
    .X(_0040_));
 sky130_fd_sc_hd__nor2_2 _0910_ (.A(_0090_),
    .B(_0462_),
    .Y(_0465_));
 sky130_fd_sc_hd__mux2_1 _0911_ (.A0(net81),
    .A1(net40),
    .S(_0465_),
    .X(_0041_));
 sky130_fd_sc_hd__mux2_1 _0912_ (.A0(net93),
    .A1(net37),
    .S(_0465_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _0913_ (.A0(net75),
    .A1(net35),
    .S(_0465_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _0914_ (.A0(net82),
    .A1(net32),
    .S(_0465_),
    .X(_0044_));
 sky130_fd_sc_hd__nor2_2 _0915_ (.A(_0460_),
    .B(_0462_),
    .Y(_0466_));
 sky130_fd_sc_hd__mux2_1 _0916_ (.A0(net85),
    .A1(net39),
    .S(_0466_),
    .X(_0045_));
 sky130_fd_sc_hd__mux2_1 _0917_ (.A0(net88),
    .A1(net37),
    .S(_0466_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _0918_ (.A0(net95),
    .A1(net35),
    .S(_0466_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _0919_ (.A0(net76),
    .A1(net32),
    .S(_0466_),
    .X(_0048_));
 sky130_fd_sc_hd__nand2b_2 _0920_ (.A_N(\counter[3] ),
    .B(\counter[2] ),
    .Y(_0467_));
 sky130_fd_sc_hd__nand3b_4 _0921_ (.A_N(\counter[3] ),
    .B(_0456_),
    .C(\counter[2] ),
    .Y(_0468_));
 sky130_fd_sc_hd__mux2_1 _0922_ (.A0(net39),
    .A1(net129),
    .S(_0468_),
    .X(_0049_));
 sky130_fd_sc_hd__mux2_1 _0923_ (.A0(net37),
    .A1(net124),
    .S(_0468_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _0924_ (.A0(net35),
    .A1(net111),
    .S(_0468_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _0925_ (.A0(net32),
    .A1(net112),
    .S(_0468_),
    .X(_0052_));
 sky130_fd_sc_hd__nor2_2 _0926_ (.A(_0089_),
    .B(_0467_),
    .Y(_0469_));
 sky130_fd_sc_hd__mux2_1 _0927_ (.A0(net96),
    .A1(net39),
    .S(_0469_),
    .X(_0053_));
 sky130_fd_sc_hd__mux2_1 _0928_ (.A0(net97),
    .A1(net7),
    .S(_0469_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _0929_ (.A0(net113),
    .A1(net36),
    .S(_0469_),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _0930_ (.A0(net83),
    .A1(net32),
    .S(_0469_),
    .X(_0056_));
 sky130_fd_sc_hd__nor2_2 _0931_ (.A(_0090_),
    .B(_0467_),
    .Y(_0470_));
 sky130_fd_sc_hd__mux2_1 _0932_ (.A0(net72),
    .A1(net40),
    .S(_0470_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _0933_ (.A0(net78),
    .A1(net7),
    .S(_0470_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _0934_ (.A0(net86),
    .A1(net35),
    .S(_0470_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _0935_ (.A0(net127),
    .A1(net32),
    .S(_0470_),
    .X(_0060_));
 sky130_fd_sc_hd__nor2_1 _0936_ (.A(_0460_),
    .B(_0467_),
    .Y(_0471_));
 sky130_fd_sc_hd__mux2_1 _0937_ (.A0(net123),
    .A1(net41),
    .S(_0471_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _0938_ (.A0(net79),
    .A1(net7),
    .S(_0471_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _0939_ (.A0(net107),
    .A1(net8),
    .S(_0471_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _0940_ (.A0(net122),
    .A1(net34),
    .S(_0471_),
    .X(_0064_));
 sky130_fd_sc_hd__or2_2 _0941_ (.A(\counter[2] ),
    .B(\counter[3] ),
    .X(_0472_));
 sky130_fd_sc_hd__or3b_2 _0942_ (.A(\counter[2] ),
    .B(\counter[3] ),
    .C_N(_0456_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_1 _0943_ (.A0(net39),
    .A1(net130),
    .S(_0473_),
    .X(_0065_));
 sky130_fd_sc_hd__mux2_1 _0944_ (.A0(net37),
    .A1(net126),
    .S(_0473_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _0945_ (.A0(net8),
    .A1(net108),
    .S(_0473_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _0946_ (.A0(net32),
    .A1(net105),
    .S(_0473_),
    .X(_0068_));
 sky130_fd_sc_hd__nor2_2 _0947_ (.A(_0089_),
    .B(_0472_),
    .Y(_0474_));
 sky130_fd_sc_hd__mux2_1 _0948_ (.A0(net103),
    .A1(net39),
    .S(_0474_),
    .X(_0069_));
 sky130_fd_sc_hd__mux2_1 _0949_ (.A0(net74),
    .A1(net38),
    .S(_0474_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _0950_ (.A0(net99),
    .A1(net35),
    .S(_0474_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _0951_ (.A0(net73),
    .A1(net32),
    .S(_0474_),
    .X(_0072_));
 sky130_fd_sc_hd__nor2_2 _0952_ (.A(_0090_),
    .B(_0472_),
    .Y(_0475_));
 sky130_fd_sc_hd__mux2_1 _0953_ (.A0(net131),
    .A1(net41),
    .S(_0475_),
    .X(_0073_));
 sky130_fd_sc_hd__mux2_1 _0954_ (.A0(net89),
    .A1(net7),
    .S(_0475_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _0955_ (.A0(net117),
    .A1(net8),
    .S(_0475_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _0956_ (.A0(net125),
    .A1(net34),
    .S(_0475_),
    .X(_0076_));
 sky130_fd_sc_hd__nor2_2 _0957_ (.A(_0460_),
    .B(_0472_),
    .Y(_0476_));
 sky130_fd_sc_hd__mux2_1 _0958_ (.A0(net102),
    .A1(net39),
    .S(_0476_),
    .X(_0077_));
 sky130_fd_sc_hd__mux2_1 _0959_ (.A0(net92),
    .A1(net38),
    .S(_0476_),
    .X(_0078_));
 sky130_fd_sc_hd__mux2_1 _0960_ (.A0(net132),
    .A1(net36),
    .S(_0476_),
    .X(_0079_));
 sky130_fd_sc_hd__mux2_1 _0961_ (.A0(net98),
    .A1(net33),
    .S(_0476_),
    .X(_0080_));
 sky130_fd_sc_hd__mux2_1 _0962_ (.A0(net42),
    .A1(\start_seg[0] ),
    .S(_0448_),
    .X(_0081_));
 sky130_fd_sc_hd__mux2_1 _0963_ (.A0(net3),
    .A1(\start_seg[1] ),
    .S(_0448_),
    .X(_0082_));
 sky130_fd_sc_hd__a21o_1 _0964_ (.A1(\start_seg[2] ),
    .A2(_0448_),
    .B1(_0451_),
    .X(_0083_));
 sky130_fd_sc_hd__mux2_1 _0965_ (.A0(net5),
    .A1(\start_seg[3] ),
    .S(_0448_),
    .X(_0084_));
 sky130_fd_sc_hd__dfrtp_1 _0966_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0012_),
    .RESET_B(net53),
    .Q(mode_dec));
 sky130_fd_sc_hd__dfrtp_1 _0967_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0013_),
    .RESET_B(net49),
    .Q(\curr_seg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _0968_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0014_),
    .RESET_B(net51),
    .Q(\curr_seg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _0969_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0015_),
    .RESET_B(net49),
    .Q(\curr_seg[2] ));
 sky130_fd_sc_hd__dfrtp_1 _0970_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0016_),
    .RESET_B(net52),
    .Q(\curr_seg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _0971_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0017_),
    .RESET_B(net44),
    .Q(\key_bytes[0][4] ));
 sky130_fd_sc_hd__dfrtp_1 _0972_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0018_),
    .RESET_B(net47),
    .Q(\key_bytes[0][5] ));
 sky130_fd_sc_hd__dfrtp_1 _0973_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0019_),
    .RESET_B(net44),
    .Q(\key_bytes[0][6] ));
 sky130_fd_sc_hd__dfrtp_1 _0974_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0020_),
    .RESET_B(net47),
    .Q(\key_bytes[0][7] ));
 sky130_fd_sc_hd__dfrtp_1 _0975_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0021_),
    .RESET_B(net46),
    .Q(\key_bytes[1][4] ));
 sky130_fd_sc_hd__dfrtp_1 _0976_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0022_),
    .RESET_B(net43),
    .Q(\key_bytes[1][5] ));
 sky130_fd_sc_hd__dfrtp_1 _0977_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0023_),
    .RESET_B(net43),
    .Q(\key_bytes[1][6] ));
 sky130_fd_sc_hd__dfrtp_1 _0978_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0024_),
    .RESET_B(net46),
    .Q(\key_bytes[1][7] ));
 sky130_fd_sc_hd__dfrtp_1 _0979_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0025_),
    .RESET_B(net50),
    .Q(\key_bytes[2][4] ));
 sky130_fd_sc_hd__dfrtp_1 _0980_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0026_),
    .RESET_B(net49),
    .Q(\key_bytes[2][5] ));
 sky130_fd_sc_hd__dfrtp_1 _0981_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0027_),
    .RESET_B(net49),
    .Q(\key_bytes[2][6] ));
 sky130_fd_sc_hd__dfrtp_1 _0982_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0028_),
    .RESET_B(net50),
    .Q(\key_bytes[2][7] ));
 sky130_fd_sc_hd__dfrtp_1 _0983_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0029_),
    .RESET_B(net50),
    .Q(\key_bytes[3][4] ));
 sky130_fd_sc_hd__dfrtp_1 _0984_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0030_),
    .RESET_B(net50),
    .Q(\key_bytes[3][5] ));
 sky130_fd_sc_hd__dfrtp_1 _0985_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0031_),
    .RESET_B(net49),
    .Q(\key_bytes[3][6] ));
 sky130_fd_sc_hd__dfrtp_1 _0986_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0032_),
    .RESET_B(net50),
    .Q(\key_bytes[3][7] ));
 sky130_fd_sc_hd__dfrtp_1 _0987_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0033_),
    .RESET_B(net46),
    .Q(\key_bytes[4][4] ));
 sky130_fd_sc_hd__dfrtp_1 _0988_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0034_),
    .RESET_B(net49),
    .Q(\key_bytes[4][5] ));
 sky130_fd_sc_hd__dfrtp_1 _0989_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0035_),
    .RESET_B(net49),
    .Q(\key_bytes[4][6] ));
 sky130_fd_sc_hd__dfrtp_1 _0990_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0036_),
    .RESET_B(net46),
    .Q(\key_bytes[4][7] ));
 sky130_fd_sc_hd__dfrtp_1 _0991_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0037_),
    .RESET_B(net43),
    .Q(\key_bytes[5][4] ));
 sky130_fd_sc_hd__dfrtp_1 _0992_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0038_),
    .RESET_B(net43),
    .Q(\key_bytes[5][5] ));
 sky130_fd_sc_hd__dfrtp_1 _0993_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0039_),
    .RESET_B(net43),
    .Q(\key_bytes[5][6] ));
 sky130_fd_sc_hd__dfrtp_1 _0994_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0040_),
    .RESET_B(net46),
    .Q(\key_bytes[5][7] ));
 sky130_fd_sc_hd__dfrtp_1 _0995_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0041_),
    .RESET_B(net47),
    .Q(\key_bytes[6][4] ));
 sky130_fd_sc_hd__dfrtp_1 _0996_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0042_),
    .RESET_B(net44),
    .Q(\key_bytes[6][5] ));
 sky130_fd_sc_hd__dfrtp_1 _0997_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0043_),
    .RESET_B(net43),
    .Q(\key_bytes[6][6] ));
 sky130_fd_sc_hd__dfrtp_1 _0998_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0044_),
    .RESET_B(net47),
    .Q(\key_bytes[6][7] ));
 sky130_fd_sc_hd__dfrtp_1 _0999_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0045_),
    .RESET_B(net44),
    .Q(\key_bytes[7][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1000_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0046_),
    .RESET_B(net44),
    .Q(\key_bytes[7][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1001_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0047_),
    .RESET_B(net43),
    .Q(\key_bytes[7][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1002_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0048_),
    .RESET_B(net46),
    .Q(\key_bytes[7][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1003_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0049_),
    .RESET_B(net44),
    .Q(\key_bytes[8][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1004_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0050_),
    .RESET_B(net43),
    .Q(\key_bytes[8][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1005_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0051_),
    .RESET_B(net43),
    .Q(\key_bytes[8][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1006_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0052_),
    .RESET_B(net46),
    .Q(\key_bytes[8][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1007_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0053_),
    .RESET_B(net45),
    .Q(\key_bytes[9][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1008_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0054_),
    .RESET_B(net49),
    .Q(\key_bytes[9][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1009_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0055_),
    .RESET_B(net49),
    .Q(\key_bytes[9][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1010_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0056_),
    .RESET_B(net46),
    .Q(\key_bytes[9][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1011_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0057_),
    .RESET_B(net47),
    .Q(\key_bytes[10][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1012_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0058_),
    .RESET_B(net49),
    .Q(\key_bytes[10][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1013_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0059_),
    .RESET_B(net45),
    .Q(\key_bytes[10][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1014_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0060_),
    .RESET_B(net46),
    .Q(\key_bytes[10][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1015_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0061_),
    .RESET_B(net50),
    .Q(\key_bytes[11][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1016_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0062_),
    .RESET_B(net50),
    .Q(\key_bytes[11][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1017_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0063_),
    .RESET_B(net50),
    .Q(\key_bytes[11][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1018_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0064_),
    .RESET_B(net50),
    .Q(\key_bytes[11][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1019_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0065_),
    .RESET_B(net44),
    .Q(\key_bytes[12][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1020_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0066_),
    .RESET_B(net43),
    .Q(\key_bytes[12][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1021_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0067_),
    .RESET_B(net52),
    .Q(\key_bytes[12][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1022_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0068_),
    .RESET_B(net46),
    .Q(\key_bytes[12][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1023_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0069_),
    .RESET_B(net45),
    .Q(\key_bytes[13][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1024_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0070_),
    .RESET_B(net45),
    .Q(\key_bytes[13][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1025_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0071_),
    .RESET_B(net45),
    .Q(\key_bytes[13][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1026_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0072_),
    .RESET_B(net47),
    .Q(\key_bytes[13][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1027_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0073_),
    .RESET_B(net50),
    .Q(\key_bytes[14][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1028_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0074_),
    .RESET_B(net52),
    .Q(\key_bytes[14][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1029_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0075_),
    .RESET_B(net51),
    .Q(\key_bytes[14][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1030_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0076_),
    .RESET_B(net51),
    .Q(\key_bytes[14][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1031_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0077_),
    .RESET_B(net44),
    .Q(\key_bytes[15][4] ));
 sky130_fd_sc_hd__dfrtp_1 _1032_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0078_),
    .RESET_B(net44),
    .Q(\key_bytes[15][5] ));
 sky130_fd_sc_hd__dfrtp_1 _1033_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0079_),
    .RESET_B(net44),
    .Q(\key_bytes[15][6] ));
 sky130_fd_sc_hd__dfrtp_1 _1034_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0080_),
    .RESET_B(net47),
    .Q(\key_bytes[15][7] ));
 sky130_fd_sc_hd__dfrtp_1 _1035_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0000_),
    .RESET_B(net51),
    .Q(\counter[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1036_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0001_),
    .RESET_B(net51),
    .Q(\counter[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1037_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0002_),
    .RESET_B(net51),
    .Q(\counter[2] ));
 sky130_fd_sc_hd__dfrtp_4 _1038_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0003_),
    .RESET_B(net51),
    .Q(\counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1039_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0004_),
    .RESET_B(net53),
    .Q(\feistel_out_q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1040_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0005_),
    .RESET_B(net53),
    .Q(\feistel_out_q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1041_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0006_),
    .RESET_B(net48),
    .Q(\feistel_out_q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1042_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0007_),
    .RESET_B(net53),
    .Q(\feistel_out_q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1043_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0008_),
    .RESET_B(net53),
    .Q(\feistel_out_q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1044_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0009_),
    .RESET_B(net48),
    .Q(\feistel_out_q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1045_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0010_),
    .RESET_B(net48),
    .Q(\feistel_out_q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1046_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0011_),
    .RESET_B(net48),
    .Q(\feistel_out_q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1047_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0477_),
    .RESET_B(net53),
    .Q(prev_streaming));
 sky130_fd_sc_hd__dfrtp_2 _1048_ (.CLK(clknet_3_7__leaf_clk),
    .D(net70),
    .RESET_B(net53),
    .Q(out_valid));
 sky130_fd_sc_hd__dfrtp_2 _1049_ (.CLK(clknet_3_5__leaf_clk),
    .D(\sys_next_state[0] ),
    .RESET_B(net51),
    .Q(\sys_state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1050_ (.CLK(clknet_3_7__leaf_clk),
    .D(\sys_next_state[1] ),
    .RESET_B(net51),
    .Q(\sys_state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1051_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0081_),
    .RESET_B(net53),
    .Q(\start_seg[0] ));
 sky130_fd_sc_hd__dfrtp_4 _1052_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0082_),
    .RESET_B(net53),
    .Q(\start_seg[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1053_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0083_),
    .RESET_B(net1),
    .Q(\start_seg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1054_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0084_),
    .RESET_B(net47),
    .Q(\start_seg[3] ));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_62 (.LO(net62));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_63 (.LO(net63));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_64 (.LO(net64));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_65 (.LO(net65));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_66 (.LO(net66));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_67 (.LO(net67));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_68 (.LO(net68));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_69 (.LO(net69));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 ();
 sky130_fd_sc_hd__dlymetal6s2s_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__buf_1 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_4 input5 (.A(ui_in[3]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_2 input7 (.A(ui_in[5]),
    .X(net7));
 sky130_fd_sc_hd__dlymetal6s2s_1 input8 (.A(ui_in[6]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 max_cap12 (.A(_0198_),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_4 fanout13 (.A(_0170_),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(_0139_),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_2 fanout15 (.A(_0139_),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_4 fanout16 (.A(_0138_),
    .X(net16));
 sky130_fd_sc_hd__buf_1 max_cap17 (.A(_0117_),
    .X(net17));
 sky130_fd_sc_hd__buf_1 wire18 (.A(_0115_),
    .X(net18));
 sky130_fd_sc_hd__buf_1 max_cap19 (.A(_0114_),
    .X(net19));
 sky130_fd_sc_hd__buf_1 max_cap20 (.A(_0095_),
    .X(net20));
 sky130_fd_sc_hd__buf_2 fanout21 (.A(_0477_),
    .X(net21));
 sky130_fd_sc_hd__buf_2 fanout22 (.A(\sys_state[1] ),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_2 fanout23 (.A(\curr_seg[3] ),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_2 fanout24 (.A(\curr_seg[3] ),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_2 fanout25 (.A(net26),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_2 fanout26 (.A(\curr_seg[2] ),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_2 fanout27 (.A(net28),
    .X(net27));
 sky130_fd_sc_hd__buf_2 fanout28 (.A(\curr_seg[1] ),
    .X(net28));
 sky130_fd_sc_hd__clkbuf_2 fanout29 (.A(net30),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(\curr_seg[0] ),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(mode_dec),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net34),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(net9),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net36),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net8),
    .X(net36));
 sky130_fd_sc_hd__buf_2 fanout37 (.A(net38),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_4 fanout38 (.A(net7),
    .X(net38));
 sky130_fd_sc_hd__buf_2 fanout39 (.A(net40),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__buf_2 fanout41 (.A(net6),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net2),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net45),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_2 fanout45 (.A(net48),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_4 fanout46 (.A(net47),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_4 fanout47 (.A(net48),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_2 fanout48 (.A(net1),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 fanout49 (.A(net52),
    .X(net49));
 sky130_fd_sc_hd__clkbuf_4 fanout50 (.A(net51),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 fanout51 (.A(net52),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_2 fanout52 (.A(net53),
    .X(net52));
 sky130_fd_sc_hd__clkbuf_4 fanout53 (.A(net1),
    .X(net53));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_54 (.LO(net54));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload3 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload4 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__inv_8 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(prev_streaming),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\key_bytes[0][5] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\key_bytes[10][4] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\key_bytes[13][7] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\key_bytes[13][5] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\key_bytes[6][6] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\key_bytes[7][7] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\key_bytes[2][4] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\key_bytes[10][5] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\key_bytes[11][5] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\key_bytes[2][7] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\key_bytes[6][4] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\key_bytes[6][7] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\key_bytes[9][7] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\key_bytes[2][6] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\key_bytes[7][4] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\key_bytes[10][6] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\key_bytes[5][7] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\key_bytes[7][5] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\key_bytes[14][5] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\key_bytes[5][5] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\key_bytes[2][5] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\key_bytes[15][5] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\key_bytes[6][5] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\key_bytes[1][4] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\key_bytes[7][6] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\key_bytes[9][4] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\key_bytes[9][5] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\key_bytes[15][7] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\key_bytes[13][6] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\key_bytes[3][5] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\key_bytes[4][4] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\key_bytes[15][4] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\key_bytes[13][4] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\key_bytes[4][5] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\key_bytes[12][7] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\key_bytes[3][7] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\key_bytes[11][6] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\key_bytes[12][6] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\key_bytes[3][6] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\key_bytes[5][4] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\key_bytes[8][6] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\key_bytes[8][7] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\key_bytes[9][6] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\key_bytes[1][6] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\key_bytes[4][7] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\key_bytes[4][6] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\key_bytes[14][6] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\key_bytes[3][4] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\key_bytes[1][5] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\key_bytes[0][4] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\key_bytes[5][6] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\key_bytes[11][7] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\key_bytes[11][4] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\key_bytes[8][5] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\key_bytes[14][7] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\key_bytes[12][5] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\key_bytes[10][7] ),
    .X(net127));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\key_bytes[1][7] ),
    .X(net128));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\key_bytes[8][4] ),
    .X(net129));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\key_bytes[12][4] ),
    .X(net130));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\key_bytes[14][4] ),
    .X(net131));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\key_bytes[15][6] ),
    .X(net132));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\key_bytes[0][6] ),
    .X(net133));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\counter[0] ),
    .X(net134));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_127 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_164 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_180 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_159 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_297 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_77 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_3_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_112 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_191 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_199 ();
 sky130_fd_sc_hd__fill_2 FILLER_5_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_78 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_161 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_261 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_7_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_80 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_86 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_208 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_139 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_172 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_235 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_10_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_184 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_92 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_96 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_141 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_238 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_299 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_173 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_245 ();
 sky130_fd_sc_hd__fill_2 FILLER_13_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_128 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_138 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_14_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_86 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_191 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_222 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_89 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_17_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_18_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_240 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_261 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_110 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_148 ();
 sky130_fd_sc_hd__decap_8 FILLER_20_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_234 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_270 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_132 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_194 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_70 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_205 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_127 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_204 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_256 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_283 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_291 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_35 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_45 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_54 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_74 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_86 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_131 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_275 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_64 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_177 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_266 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_135 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_27_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_49 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_163 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_188 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_207 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_215 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_156 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_201 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_60 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_176 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_30_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_263 ();
 sky130_fd_sc_hd__decap_3 FILLER_30_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_133 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_146 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_255 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_267 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_206 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_210 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_32_249 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_284 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_33_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_123 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_168 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_236 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_294 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_151 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_278 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_36_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_217 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_236 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_250 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_166 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_189 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_148 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_162 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_273 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_331 ();
 assign uio_oe[0] = net54;
 assign uio_oe[1] = net55;
 assign uio_oe[2] = net56;
 assign uio_oe[3] = net57;
 assign uio_oe[4] = net58;
 assign uio_oe[5] = net59;
 assign uio_oe[6] = net60;
 assign uio_oe[7] = net61;
 assign uio_out[0] = net62;
 assign uio_out[1] = net63;
 assign uio_out[2] = net64;
 assign uio_out[3] = net65;
 assign uio_out[4] = net66;
 assign uio_out[5] = net67;
 assign uio_out[6] = net68;
 assign uio_out[7] = net69;
endmodule
