module tt_um_Samcooper01 (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire \counter[0] ;
 wire \counter[1] ;
 wire \counter[2] ;
 wire \counter[3] ;
 wire \counter[4] ;
 wire \curr_seg[0] ;
 wire \curr_seg[1] ;
 wire \curr_seg[2] ;
 wire \curr_seg[3] ;
 wire \full_key[100] ;
 wire \full_key[101] ;
 wire \full_key[102] ;
 wire \full_key[103] ;
 wire \full_key[108] ;
 wire \full_key[109] ;
 wire \full_key[110] ;
 wire \full_key[111] ;
 wire \full_key[116] ;
 wire \full_key[117] ;
 wire \full_key[118] ;
 wire \full_key[119] ;
 wire \full_key[124] ;
 wire \full_key[125] ;
 wire \full_key[126] ;
 wire \full_key[127] ;
 wire \full_key[12] ;
 wire \full_key[13] ;
 wire \full_key[14] ;
 wire \full_key[15] ;
 wire \full_key[20] ;
 wire \full_key[21] ;
 wire \full_key[22] ;
 wire \full_key[23] ;
 wire \full_key[28] ;
 wire \full_key[29] ;
 wire \full_key[30] ;
 wire \full_key[31] ;
 wire \full_key[36] ;
 wire \full_key[37] ;
 wire \full_key[38] ;
 wire \full_key[39] ;
 wire \full_key[44] ;
 wire \full_key[45] ;
 wire \full_key[46] ;
 wire \full_key[47] ;
 wire \full_key[4] ;
 wire \full_key[52] ;
 wire \full_key[53] ;
 wire \full_key[54] ;
 wire \full_key[55] ;
 wire \full_key[5] ;
 wire \full_key[60] ;
 wire \full_key[61] ;
 wire \full_key[62] ;
 wire \full_key[63] ;
 wire \full_key[68] ;
 wire \full_key[69] ;
 wire \full_key[6] ;
 wire \full_key[70] ;
 wire \full_key[71] ;
 wire \full_key[76] ;
 wire \full_key[77] ;
 wire \full_key[78] ;
 wire \full_key[79] ;
 wire \full_key[7] ;
 wire \full_key[84] ;
 wire \full_key[85] ;
 wire \full_key[86] ;
 wire \full_key[87] ;
 wire \full_key[92] ;
 wire \full_key[93] ;
 wire \full_key[94] ;
 wire \full_key[95] ;
 wire mode_dec;
 wire \start_seg[0] ;
 wire \start_seg[1] ;
 wire \start_seg[2] ;
 wire \start_seg[3] ;
 wire \sys_next_state[0] ;
 wire \sys_next_state[1] ;
 wire \sys_state[0] ;
 wire \sys_state[1] ;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire clknet_0_clk;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;

 sky130_fd_sc_hd__inv_2 _0529_ (.A(net2),
    .Y(_0078_));
 sky130_fd_sc_hd__inv_2 _0530_ (.A(net23),
    .Y(_0079_));
 sky130_fd_sc_hd__inv_2 _0531_ (.A(\curr_seg[3] ),
    .Y(_0080_));
 sky130_fd_sc_hd__inv_2 _0532_ (.A(net3),
    .Y(_0081_));
 sky130_fd_sc_hd__inv_2 _0533_ (.A(\start_seg[1] ),
    .Y(_0082_));
 sky130_fd_sc_hd__inv_2 _0534_ (.A(mode_dec),
    .Y(_0083_));
 sky130_fd_sc_hd__inv_2 _0535_ (.A(net11),
    .Y(_0084_));
 sky130_fd_sc_hd__and2_1 _0536_ (.A(net20),
    .B(\sys_state[0] ),
    .X(_0085_));
 sky130_fd_sc_hd__nand2_4 _0537_ (.A(net20),
    .B(\sys_state[0] ),
    .Y(_0086_));
 sky130_fd_sc_hd__nand2_4 _0538_ (.A(net28),
    .B(net19),
    .Y(_0087_));
 sky130_fd_sc_hd__nand2_1 _0539_ (.A(net2),
    .B(net18),
    .Y(_0088_));
 sky130_fd_sc_hd__inv_2 _0540_ (.A(_0088_),
    .Y(_0089_));
 sky130_fd_sc_hd__o22a_1 _0541_ (.A1(net2),
    .A2(_0087_),
    .B1(_0088_),
    .B2(net28),
    .X(_0090_));
 sky130_fd_sc_hd__and3_1 _0542_ (.A(net20),
    .B(\sys_state[0] ),
    .C(net31),
    .X(_0091_));
 sky130_fd_sc_hd__nand2_1 _0543_ (.A(net30),
    .B(net18),
    .Y(_0092_));
 sky130_fd_sc_hd__mux4_1 _0544_ (.A0(\full_key[126] ),
    .A1(\full_key[118] ),
    .A2(\full_key[110] ),
    .A3(\full_key[102] ),
    .S0(net26),
    .S1(net24),
    .X(_0093_));
 sky130_fd_sc_hd__mux4_1 _0545_ (.A0(\full_key[94] ),
    .A1(\full_key[86] ),
    .A2(\full_key[78] ),
    .A3(\full_key[70] ),
    .S0(net27),
    .S1(net25),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _0546_ (.A0(_0093_),
    .A1(_0094_),
    .S(net23),
    .X(_0095_));
 sky130_fd_sc_hd__mux4_1 _0547_ (.A0(\full_key[30] ),
    .A1(\full_key[22] ),
    .A2(\full_key[14] ),
    .A3(\full_key[6] ),
    .S0(net27),
    .S1(net25),
    .X(_0096_));
 sky130_fd_sc_hd__mux4_1 _0548_ (.A0(\full_key[62] ),
    .A1(\full_key[54] ),
    .A2(\full_key[46] ),
    .A3(\full_key[38] ),
    .S0(net26),
    .S1(net24),
    .X(_0097_));
 sky130_fd_sc_hd__or2_1 _0549_ (.A(net23),
    .B(_0097_),
    .X(_0098_));
 sky130_fd_sc_hd__o21a_1 _0550_ (.A1(_0079_),
    .A2(_0096_),
    .B1(\curr_seg[3] ),
    .X(_0099_));
 sky130_fd_sc_hd__a22o_1 _0551_ (.A1(_0080_),
    .A2(_0095_),
    .B1(_0098_),
    .B2(_0099_),
    .X(_0100_));
 sky130_fd_sc_hd__and3_4 _0552_ (.A(net20),
    .B(\sys_state[0] ),
    .C(net46),
    .X(_0101_));
 sky130_fd_sc_hd__nand2_1 _0553_ (.A(net46),
    .B(net18),
    .Y(_0102_));
 sky130_fd_sc_hd__or3b_2 _0554_ (.A(\start_seg[2] ),
    .B(_0102_),
    .C_N(_0100_),
    .X(_0103_));
 sky130_fd_sc_hd__a21bo_1 _0555_ (.A1(_0100_),
    .A2(_0101_),
    .B1_N(\start_seg[2] ),
    .X(_0104_));
 sky130_fd_sc_hd__and2_4 _0556_ (.A(_0103_),
    .B(_0104_),
    .X(_0105_));
 sky130_fd_sc_hd__inv_2 _0557_ (.A(_0105_),
    .Y(_0106_));
 sky130_fd_sc_hd__nand2_1 _0558_ (.A(\start_seg[0] ),
    .B(\start_seg[1] ),
    .Y(_0107_));
 sky130_fd_sc_hd__a21bo_1 _0559_ (.A1(_0103_),
    .A2(_0104_),
    .B1_N(_0107_),
    .X(_0108_));
 sky130_fd_sc_hd__nand3b_2 _0560_ (.A_N(_0107_),
    .B(_0104_),
    .C(_0103_),
    .Y(_0109_));
 sky130_fd_sc_hd__nand2_4 _0561_ (.A(_0108_),
    .B(_0109_),
    .Y(_0110_));
 sky130_fd_sc_hd__and3_1 _0562_ (.A(_0091_),
    .B(_0108_),
    .C(_0109_),
    .X(_0111_));
 sky130_fd_sc_hd__a21oi_1 _0563_ (.A1(_0108_),
    .A2(_0109_),
    .B1(_0091_),
    .Y(_0112_));
 sky130_fd_sc_hd__mux4_1 _0564_ (.A0(\full_key[61] ),
    .A1(\full_key[53] ),
    .A2(\full_key[45] ),
    .A3(\full_key[37] ),
    .S0(net26),
    .S1(net24),
    .X(_0113_));
 sky130_fd_sc_hd__or2_1 _0565_ (.A(net23),
    .B(_0113_),
    .X(_0114_));
 sky130_fd_sc_hd__mux4_1 _0566_ (.A0(\full_key[29] ),
    .A1(\full_key[21] ),
    .A2(\full_key[13] ),
    .A3(\full_key[5] ),
    .S0(net27),
    .S1(net25),
    .X(_0115_));
 sky130_fd_sc_hd__o21a_1 _0567_ (.A1(_0079_),
    .A2(_0115_),
    .B1(\curr_seg[3] ),
    .X(_0116_));
 sky130_fd_sc_hd__mux4_1 _0568_ (.A0(\full_key[125] ),
    .A1(\full_key[117] ),
    .A2(\full_key[109] ),
    .A3(\full_key[101] ),
    .S0(net26),
    .S1(net24),
    .X(_0117_));
 sky130_fd_sc_hd__mux4_1 _0569_ (.A0(\full_key[93] ),
    .A1(\full_key[85] ),
    .A2(\full_key[77] ),
    .A3(\full_key[69] ),
    .S0(net26),
    .S1(net24),
    .X(_0118_));
 sky130_fd_sc_hd__mux2_1 _0570_ (.A0(_0117_),
    .A1(_0118_),
    .S(net23),
    .X(_0119_));
 sky130_fd_sc_hd__a22o_1 _0571_ (.A1(_0114_),
    .A2(_0116_),
    .B1(_0119_),
    .B2(_0080_),
    .X(_0120_));
 sky130_fd_sc_hd__or2_1 _0572_ (.A(\start_seg[0] ),
    .B(\start_seg[1] ),
    .X(_0121_));
 sky130_fd_sc_hd__nand2_1 _0573_ (.A(_0107_),
    .B(_0121_),
    .Y(_0122_));
 sky130_fd_sc_hd__nand3_1 _0574_ (.A(_0101_),
    .B(_0120_),
    .C(_0122_),
    .Y(_0123_));
 sky130_fd_sc_hd__a21o_1 _0575_ (.A1(_0101_),
    .A2(_0120_),
    .B1(_0122_),
    .X(_0124_));
 sky130_fd_sc_hd__nand2_1 _0576_ (.A(_0123_),
    .B(_0124_),
    .Y(_0125_));
 sky130_fd_sc_hd__and2_1 _0577_ (.A(_0123_),
    .B(_0124_),
    .X(_0126_));
 sky130_fd_sc_hd__nand2_1 _0578_ (.A(net32),
    .B(net18),
    .Y(_0127_));
 sky130_fd_sc_hd__and3_1 _0579_ (.A(_0123_),
    .B(_0124_),
    .C(_0127_),
    .X(_0128_));
 sky130_fd_sc_hd__a21oi_1 _0580_ (.A1(_0123_),
    .A2(_0124_),
    .B1(_0127_),
    .Y(_0129_));
 sky130_fd_sc_hd__mux4_1 _0581_ (.A0(\full_key[60] ),
    .A1(\full_key[52] ),
    .A2(\full_key[44] ),
    .A3(\full_key[36] ),
    .S0(net26),
    .S1(net24),
    .X(_0130_));
 sky130_fd_sc_hd__or2_1 _0582_ (.A(\curr_seg[2] ),
    .B(_0130_),
    .X(_0131_));
 sky130_fd_sc_hd__mux4_1 _0583_ (.A0(\full_key[28] ),
    .A1(\full_key[20] ),
    .A2(\full_key[12] ),
    .A3(\full_key[4] ),
    .S0(net27),
    .S1(net25),
    .X(_0132_));
 sky130_fd_sc_hd__o21a_1 _0584_ (.A1(_0079_),
    .A2(_0132_),
    .B1(\curr_seg[3] ),
    .X(_0133_));
 sky130_fd_sc_hd__mux4_1 _0585_ (.A0(\full_key[124] ),
    .A1(\full_key[116] ),
    .A2(\full_key[108] ),
    .A3(\full_key[100] ),
    .S0(net26),
    .S1(net24),
    .X(_0134_));
 sky130_fd_sc_hd__mux4_1 _0586_ (.A0(\full_key[92] ),
    .A1(\full_key[84] ),
    .A2(\full_key[76] ),
    .A3(\full_key[68] ),
    .S0(net26),
    .S1(net24),
    .X(_0135_));
 sky130_fd_sc_hd__mux2_1 _0587_ (.A0(_0134_),
    .A1(_0135_),
    .S(net23),
    .X(_0136_));
 sky130_fd_sc_hd__a22o_1 _0588_ (.A1(_0131_),
    .A2(_0133_),
    .B1(_0136_),
    .B2(_0080_),
    .X(_0137_));
 sky130_fd_sc_hd__and3_2 _0589_ (.A(\start_seg[0] ),
    .B(_0101_),
    .C(_0137_),
    .X(_0138_));
 sky130_fd_sc_hd__a21oi_4 _0590_ (.A1(_0101_),
    .A2(_0137_),
    .B1(\start_seg[0] ),
    .Y(_0139_));
 sky130_fd_sc_hd__or3b_1 _0591_ (.A(\start_seg[0] ),
    .B(_0102_),
    .C_N(_0137_),
    .X(_0140_));
 sky130_fd_sc_hd__a21bo_1 _0592_ (.A1(_0101_),
    .A2(_0137_),
    .B1_N(\start_seg[0] ),
    .X(_0141_));
 sky130_fd_sc_hd__nor2_1 _0593_ (.A(_0138_),
    .B(_0139_),
    .Y(_0142_));
 sky130_fd_sc_hd__or2_2 _0594_ (.A(_0138_),
    .B(_0139_),
    .X(_0143_));
 sky130_fd_sc_hd__and3_1 _0595_ (.A(net20),
    .B(\sys_state[0] ),
    .C(net34),
    .X(_0144_));
 sky130_fd_sc_hd__nand2_1 _0596_ (.A(net34),
    .B(net18),
    .Y(_0145_));
 sky130_fd_sc_hd__o21ai_2 _0597_ (.A1(_0138_),
    .A2(_0139_),
    .B1(_0144_),
    .Y(_0146_));
 sky130_fd_sc_hd__o21ba_1 _0598_ (.A1(_0128_),
    .A2(_0146_),
    .B1_N(_0129_),
    .X(_0147_));
 sky130_fd_sc_hd__or3_1 _0599_ (.A(_0111_),
    .B(_0112_),
    .C(_0147_),
    .X(_0148_));
 sky130_fd_sc_hd__o21ba_1 _0600_ (.A1(_0112_),
    .A2(_0147_),
    .B1_N(_0111_),
    .X(_0149_));
 sky130_fd_sc_hd__nand2_1 _0601_ (.A(net5),
    .B(net19),
    .Y(_0150_));
 sky130_fd_sc_hd__o22a_1 _0602_ (.A1(net5),
    .A2(_0087_),
    .B1(_0150_),
    .B2(net9),
    .X(_0151_));
 sky130_fd_sc_hd__mux2_1 _0603_ (.A0(net30),
    .A1(_0092_),
    .S(_0151_),
    .X(_0152_));
 sky130_fd_sc_hd__mux4_1 _0604_ (.A0(\full_key[63] ),
    .A1(\full_key[55] ),
    .A2(\full_key[47] ),
    .A3(\full_key[39] ),
    .S0(net26),
    .S1(net24),
    .X(_0153_));
 sky130_fd_sc_hd__or2_1 _0605_ (.A(net23),
    .B(_0153_),
    .X(_0154_));
 sky130_fd_sc_hd__mux4_1 _0606_ (.A0(\full_key[31] ),
    .A1(\full_key[23] ),
    .A2(\full_key[15] ),
    .A3(\full_key[7] ),
    .S0(net27),
    .S1(net25),
    .X(_0155_));
 sky130_fd_sc_hd__o21a_1 _0607_ (.A1(_0079_),
    .A2(_0155_),
    .B1(\curr_seg[3] ),
    .X(_0156_));
 sky130_fd_sc_hd__mux4_1 _0608_ (.A0(\full_key[127] ),
    .A1(\full_key[119] ),
    .A2(\full_key[111] ),
    .A3(\full_key[103] ),
    .S0(net26),
    .S1(net24),
    .X(_0157_));
 sky130_fd_sc_hd__mux4_1 _0609_ (.A0(\full_key[95] ),
    .A1(\full_key[87] ),
    .A2(\full_key[79] ),
    .A3(\full_key[71] ),
    .S0(net27),
    .S1(net25),
    .X(_0158_));
 sky130_fd_sc_hd__mux2_1 _0610_ (.A0(_0157_),
    .A1(_0158_),
    .S(net23),
    .X(_0159_));
 sky130_fd_sc_hd__a22o_1 _0611_ (.A1(_0154_),
    .A2(_0156_),
    .B1(_0159_),
    .B2(_0080_),
    .X(_0160_));
 sky130_fd_sc_hd__nand2_2 _0612_ (.A(_0101_),
    .B(_0160_),
    .Y(_0161_));
 sky130_fd_sc_hd__xor2_4 _0613_ (.A(\start_seg[3] ),
    .B(_0161_),
    .X(_0162_));
 sky130_fd_sc_hd__inv_2 _0614_ (.A(_0162_),
    .Y(_0163_));
 sky130_fd_sc_hd__a21oi_1 _0615_ (.A1(\start_seg[0] ),
    .A2(\start_seg[1] ),
    .B1(\start_seg[2] ),
    .Y(_0164_));
 sky130_fd_sc_hd__xnor2_1 _0616_ (.A(_0162_),
    .B(_0164_),
    .Y(_0165_));
 sky130_fd_sc_hd__xnor2_1 _0617_ (.A(_0152_),
    .B(_0165_),
    .Y(_0166_));
 sky130_fd_sc_hd__xnor2_2 _0618_ (.A(_0149_),
    .B(_0166_),
    .Y(_0167_));
 sky130_fd_sc_hd__xnor2_2 _0619_ (.A(_0090_),
    .B(_0167_),
    .Y(_0168_));
 sky130_fd_sc_hd__o21ai_1 _0620_ (.A1(_0111_),
    .A2(_0112_),
    .B1(_0147_),
    .Y(_0169_));
 sky130_fd_sc_hd__nand2_2 _0621_ (.A(net4),
    .B(net18),
    .Y(_0170_));
 sky130_fd_sc_hd__o22ai_1 _0622_ (.A1(net4),
    .A2(_0127_),
    .B1(_0170_),
    .B2(net32),
    .Y(_0171_));
 sky130_fd_sc_hd__a21o_1 _0623_ (.A1(_0148_),
    .A2(_0169_),
    .B1(_0171_),
    .X(_0172_));
 sky130_fd_sc_hd__nand3_1 _0624_ (.A(_0148_),
    .B(_0169_),
    .C(_0171_),
    .Y(_0173_));
 sky130_fd_sc_hd__and2_1 _0625_ (.A(_0172_),
    .B(_0173_),
    .X(_0174_));
 sky130_fd_sc_hd__a21o_1 _0626_ (.A1(_0172_),
    .A2(_0173_),
    .B1(_0106_),
    .X(_0175_));
 sky130_fd_sc_hd__or3b_2 _0627_ (.A(\start_seg[1] ),
    .B(_0102_),
    .C_N(_0120_),
    .X(_0176_));
 sky130_fd_sc_hd__a21o_1 _0628_ (.A1(_0101_),
    .A2(_0120_),
    .B1(_0082_),
    .X(_0177_));
 sky130_fd_sc_hd__nand2_4 _0629_ (.A(_0176_),
    .B(_0177_),
    .Y(_0178_));
 sky130_fd_sc_hd__and2_1 _0630_ (.A(_0176_),
    .B(_0177_),
    .X(_0179_));
 sky130_fd_sc_hd__nor2_1 _0631_ (.A(_0081_),
    .B(_0086_),
    .Y(_0180_));
 sky130_fd_sc_hd__nand2_1 _0632_ (.A(net3),
    .B(net18),
    .Y(_0181_));
 sky130_fd_sc_hd__or4_1 _0633_ (.A(net3),
    .B(_0138_),
    .C(_0139_),
    .D(_0145_),
    .X(_0182_));
 sky130_fd_sc_hd__o31ai_2 _0634_ (.A1(_0138_),
    .A2(_0139_),
    .A3(_0145_),
    .B1(_0180_),
    .Y(_0183_));
 sky130_fd_sc_hd__a211o_1 _0635_ (.A1(_0182_),
    .A2(_0183_),
    .B1(_0128_),
    .C1(_0129_),
    .X(_0184_));
 sky130_fd_sc_hd__o211ai_2 _0636_ (.A1(_0128_),
    .A2(_0129_),
    .B1(_0182_),
    .C1(_0183_),
    .Y(_0185_));
 sky130_fd_sc_hd__and2_1 _0637_ (.A(_0184_),
    .B(_0185_),
    .X(_0186_));
 sky130_fd_sc_hd__and3_1 _0638_ (.A(_0178_),
    .B(_0184_),
    .C(_0185_),
    .X(_0187_));
 sky130_fd_sc_hd__a21oi_1 _0639_ (.A1(_0184_),
    .A2(_0185_),
    .B1(_0178_),
    .Y(_0188_));
 sky130_fd_sc_hd__or3_2 _0640_ (.A(_0138_),
    .B(_0139_),
    .C(_0144_),
    .X(_0189_));
 sky130_fd_sc_hd__a21bo_1 _0641_ (.A1(_0146_),
    .A2(_0189_),
    .B1_N(_0090_),
    .X(_0190_));
 sky130_fd_sc_hd__nand3b_1 _0642_ (.A_N(_0090_),
    .B(_0146_),
    .C(_0189_),
    .Y(_0191_));
 sky130_fd_sc_hd__nand3_1 _0643_ (.A(net14),
    .B(_0190_),
    .C(_0191_),
    .Y(_0192_));
 sky130_fd_sc_hd__o21ba_1 _0644_ (.A1(_0188_),
    .A2(_0192_),
    .B1_N(_0187_),
    .X(_0193_));
 sky130_fd_sc_hd__nand3_1 _0645_ (.A(_0106_),
    .B(_0172_),
    .C(_0173_),
    .Y(_0194_));
 sky130_fd_sc_hd__mux2_2 _0646_ (.A0(_0175_),
    .A1(_0194_),
    .S(_0193_),
    .X(_0195_));
 sky130_fd_sc_hd__xnor2_2 _0647_ (.A(\start_seg[2] ),
    .B(_0162_),
    .Y(_0196_));
 sky130_fd_sc_hd__xnor2_2 _0648_ (.A(_0087_),
    .B(_0196_),
    .Y(_0197_));
 sky130_fd_sc_hd__xor2_1 _0649_ (.A(_0167_),
    .B(_0197_),
    .X(_0198_));
 sky130_fd_sc_hd__xnor2_1 _0650_ (.A(_0195_),
    .B(_0198_),
    .Y(_0199_));
 sky130_fd_sc_hd__xor2_2 _0651_ (.A(_0105_),
    .B(_0121_),
    .X(_0200_));
 sky130_fd_sc_hd__xnor2_1 _0652_ (.A(_0091_),
    .B(_0186_),
    .Y(_0201_));
 sky130_fd_sc_hd__xnor2_1 _0653_ (.A(_0193_),
    .B(_0201_),
    .Y(_0202_));
 sky130_fd_sc_hd__a21o_1 _0654_ (.A1(_0175_),
    .A2(_0194_),
    .B1(_0202_),
    .X(_0203_));
 sky130_fd_sc_hd__nand3_2 _0655_ (.A(_0175_),
    .B(_0194_),
    .C(_0202_),
    .Y(_0204_));
 sky130_fd_sc_hd__nand2_1 _0656_ (.A(_0203_),
    .B(_0204_),
    .Y(_0205_));
 sky130_fd_sc_hd__nand3b_1 _0657_ (.A_N(_0200_),
    .B(_0203_),
    .C(_0204_),
    .Y(_0206_));
 sky130_fd_sc_hd__nand4_1 _0658_ (.A(_0127_),
    .B(net12),
    .C(_0190_),
    .D(_0191_),
    .Y(_0207_));
 sky130_fd_sc_hd__a31o_1 _0659_ (.A1(net12),
    .A2(_0190_),
    .A3(_0191_),
    .B1(_0127_),
    .X(_0208_));
 sky130_fd_sc_hd__or4bb_1 _0660_ (.A(_0187_),
    .B(_0188_),
    .C_N(_0207_),
    .D_N(_0208_),
    .X(_0209_));
 sky130_fd_sc_hd__a2bb2o_1 _0661_ (.A1_N(_0187_),
    .A2_N(_0188_),
    .B1(_0207_),
    .B2(_0208_),
    .X(_0210_));
 sky130_fd_sc_hd__nand2_1 _0662_ (.A(_0209_),
    .B(_0210_),
    .Y(_0211_));
 sky130_fd_sc_hd__a21oi_1 _0663_ (.A1(_0209_),
    .A2(_0210_),
    .B1(net15),
    .Y(_0212_));
 sky130_fd_sc_hd__and3_1 _0664_ (.A(net15),
    .B(_0209_),
    .C(_0210_),
    .X(_0213_));
 sky130_fd_sc_hd__o211a_1 _0665_ (.A1(_0126_),
    .A2(_0211_),
    .B1(_0168_),
    .C1(net12),
    .X(_0214_));
 sky130_fd_sc_hd__or2_1 _0666_ (.A(_0212_),
    .B(_0214_),
    .X(_0215_));
 sky130_fd_sc_hd__a21bo_1 _0667_ (.A1(_0203_),
    .A2(_0204_),
    .B1_N(_0200_),
    .X(_0216_));
 sky130_fd_sc_hd__nand3_1 _0668_ (.A(_0206_),
    .B(_0215_),
    .C(_0216_),
    .Y(_0217_));
 sky130_fd_sc_hd__a21boi_1 _0669_ (.A1(_0215_),
    .A2(_0216_),
    .B1_N(_0206_),
    .Y(_0218_));
 sky130_fd_sc_hd__nand2_1 _0670_ (.A(\start_seg[2] ),
    .B(_0121_),
    .Y(_0219_));
 sky130_fd_sc_hd__xor2_2 _0671_ (.A(_0162_),
    .B(_0219_),
    .X(_0220_));
 sky130_fd_sc_hd__xor2_1 _0672_ (.A(_0167_),
    .B(_0220_),
    .X(_0221_));
 sky130_fd_sc_hd__and3_1 _0673_ (.A(_0203_),
    .B(_0204_),
    .C(_0221_),
    .X(_0222_));
 sky130_fd_sc_hd__a21oi_1 _0674_ (.A1(_0203_),
    .A2(_0204_),
    .B1(_0221_),
    .Y(_0223_));
 sky130_fd_sc_hd__nor2_1 _0675_ (.A(_0222_),
    .B(_0223_),
    .Y(_0224_));
 sky130_fd_sc_hd__xor2_1 _0676_ (.A(_0218_),
    .B(_0224_),
    .X(_0225_));
 sky130_fd_sc_hd__or3_1 _0677_ (.A(_0199_),
    .B(_0222_),
    .C(_0223_),
    .X(_0226_));
 sky130_fd_sc_hd__o21ai_1 _0678_ (.A1(_0222_),
    .A2(_0223_),
    .B1(_0199_),
    .Y(_0227_));
 sky130_fd_sc_hd__and3_1 _0679_ (.A(_0218_),
    .B(_0226_),
    .C(_0227_),
    .X(_0228_));
 sky130_fd_sc_hd__a21oi_1 _0680_ (.A1(_0226_),
    .A2(_0227_),
    .B1(_0218_),
    .Y(_0229_));
 sky130_fd_sc_hd__nor2_1 _0681_ (.A(_0228_),
    .B(_0229_),
    .Y(_0230_));
 sky130_fd_sc_hd__xnor2_2 _0682_ (.A(_0082_),
    .B(_0105_),
    .Y(_0231_));
 sky130_fd_sc_hd__inv_2 _0683_ (.A(_0231_),
    .Y(_0232_));
 sky130_fd_sc_hd__and2_1 _0684_ (.A(net14),
    .B(_0168_),
    .X(_0233_));
 sky130_fd_sc_hd__o21ai_1 _0685_ (.A1(_0212_),
    .A2(_0213_),
    .B1(_0186_),
    .Y(_0234_));
 sky130_fd_sc_hd__or3_1 _0686_ (.A(_0186_),
    .B(_0212_),
    .C(_0213_),
    .X(_0235_));
 sky130_fd_sc_hd__a21o_1 _0687_ (.A1(_0234_),
    .A2(_0235_),
    .B1(_0233_),
    .X(_0236_));
 sky130_fd_sc_hd__nand3_1 _0688_ (.A(_0233_),
    .B(_0234_),
    .C(_0235_),
    .Y(_0237_));
 sky130_fd_sc_hd__nand2_1 _0689_ (.A(_0236_),
    .B(_0237_),
    .Y(_0238_));
 sky130_fd_sc_hd__inv_2 _0690_ (.A(_0238_),
    .Y(_0239_));
 sky130_fd_sc_hd__and3_1 _0691_ (.A(_0178_),
    .B(_0236_),
    .C(_0237_),
    .X(_0240_));
 sky130_fd_sc_hd__nand3_1 _0692_ (.A(_0178_),
    .B(_0236_),
    .C(_0237_),
    .Y(_0241_));
 sky130_fd_sc_hd__a21o_1 _0693_ (.A1(_0236_),
    .A2(_0237_),
    .B1(_0178_),
    .X(_0242_));
 sky130_fd_sc_hd__xnor2_1 _0694_ (.A(_0145_),
    .B(_0197_),
    .Y(_0243_));
 sky130_fd_sc_hd__xnor2_2 _0695_ (.A(_0195_),
    .B(_0243_),
    .Y(_0244_));
 sky130_fd_sc_hd__or2_1 _0696_ (.A(net12),
    .B(_0244_),
    .X(_0245_));
 sky130_fd_sc_hd__o311a_1 _0697_ (.A1(net12),
    .A2(_0240_),
    .A3(_0244_),
    .B1(_0242_),
    .C1(_0231_),
    .X(_0246_));
 sky130_fd_sc_hd__a21o_1 _0698_ (.A1(_0206_),
    .A2(_0216_),
    .B1(_0215_),
    .X(_0247_));
 sky130_fd_sc_hd__xor2_1 _0699_ (.A(_0174_),
    .B(_0211_),
    .X(_0248_));
 sky130_fd_sc_hd__a21o_1 _0700_ (.A1(_0217_),
    .A2(_0247_),
    .B1(_0248_),
    .X(_0249_));
 sky130_fd_sc_hd__nand3_2 _0701_ (.A(_0217_),
    .B(_0247_),
    .C(_0248_),
    .Y(_0250_));
 sky130_fd_sc_hd__nand2_1 _0702_ (.A(_0249_),
    .B(_0250_),
    .Y(_0251_));
 sky130_fd_sc_hd__a211o_1 _0703_ (.A1(_0242_),
    .A2(_0245_),
    .B1(_0231_),
    .C1(_0240_),
    .X(_0252_));
 sky130_fd_sc_hd__a21o_1 _0704_ (.A1(_0249_),
    .A2(_0250_),
    .B1(_0252_),
    .X(_0253_));
 sky130_fd_sc_hd__nand3_1 _0705_ (.A(_0246_),
    .B(_0249_),
    .C(_0250_),
    .Y(_0254_));
 sky130_fd_sc_hd__nand2_1 _0706_ (.A(\start_seg[2] ),
    .B(\start_seg[1] ),
    .Y(_0255_));
 sky130_fd_sc_hd__xor2_2 _0707_ (.A(_0162_),
    .B(_0255_),
    .X(_0256_));
 sky130_fd_sc_hd__xor2_1 _0708_ (.A(_0225_),
    .B(_0256_),
    .X(_0257_));
 sky130_fd_sc_hd__a21o_1 _0709_ (.A1(_0253_),
    .A2(_0254_),
    .B1(_0257_),
    .X(_0258_));
 sky130_fd_sc_hd__nand3_1 _0710_ (.A(_0253_),
    .B(_0254_),
    .C(_0257_),
    .Y(_0259_));
 sky130_fd_sc_hd__and2_1 _0711_ (.A(_0258_),
    .B(_0259_),
    .X(_0260_));
 sky130_fd_sc_hd__a21o_1 _0712_ (.A1(_0258_),
    .A2(_0259_),
    .B1(_0230_),
    .X(_0261_));
 sky130_fd_sc_hd__nand3_2 _0713_ (.A(_0230_),
    .B(_0258_),
    .C(_0259_),
    .Y(_0262_));
 sky130_fd_sc_hd__nand3_1 _0714_ (.A(_0168_),
    .B(_0261_),
    .C(_0262_),
    .Y(_0263_));
 sky130_fd_sc_hd__a21o_1 _0715_ (.A1(_0261_),
    .A2(_0262_),
    .B1(_0168_),
    .X(_0264_));
 sky130_fd_sc_hd__and2_1 _0716_ (.A(_0263_),
    .B(_0264_),
    .X(_0265_));
 sky130_fd_sc_hd__a21oi_1 _0717_ (.A1(_0103_),
    .A2(_0104_),
    .B1(_0170_),
    .Y(_0266_));
 sky130_fd_sc_hd__and3_1 _0718_ (.A(_0103_),
    .B(_0104_),
    .C(_0170_),
    .X(_0267_));
 sky130_fd_sc_hd__nor2_1 _0719_ (.A(_0266_),
    .B(_0267_),
    .Y(_0268_));
 sky130_fd_sc_hd__a21oi_1 _0720_ (.A1(_0176_),
    .A2(_0177_),
    .B1(_0181_),
    .Y(_0269_));
 sky130_fd_sc_hd__and3_1 _0721_ (.A(_0176_),
    .B(_0177_),
    .C(_0181_),
    .X(_0270_));
 sky130_fd_sc_hd__or3_1 _0722_ (.A(_0088_),
    .B(_0138_),
    .C(_0139_),
    .X(_0271_));
 sky130_fd_sc_hd__o32a_1 _0723_ (.A1(_0081_),
    .A2(_0086_),
    .A3(_0179_),
    .B1(_0270_),
    .B2(_0271_),
    .X(_0272_));
 sky130_fd_sc_hd__xnor2_2 _0724_ (.A(_0268_),
    .B(_0272_),
    .Y(_0273_));
 sky130_fd_sc_hd__o22a_1 _0725_ (.A1(net3),
    .A2(_0092_),
    .B1(_0181_),
    .B2(net8),
    .X(_0274_));
 sky130_fd_sc_hd__xnor2_2 _0726_ (.A(_0273_),
    .B(_0274_),
    .Y(_0275_));
 sky130_fd_sc_hd__xor2_1 _0727_ (.A(_0273_),
    .B(_0274_),
    .X(_0276_));
 sky130_fd_sc_hd__xnor2_2 _0728_ (.A(_0110_),
    .B(_0275_),
    .Y(_0277_));
 sky130_fd_sc_hd__a32o_1 _0729_ (.A1(_0089_),
    .A2(_0140_),
    .A3(_0141_),
    .B1(net18),
    .B2(net7),
    .X(_0278_));
 sky130_fd_sc_hd__o211ai_2 _0730_ (.A1(_0138_),
    .A2(_0139_),
    .B1(net7),
    .C1(_0089_),
    .Y(_0279_));
 sky130_fd_sc_hd__a211o_1 _0731_ (.A1(_0278_),
    .A2(_0279_),
    .B1(_0269_),
    .C1(_0270_),
    .X(_0280_));
 sky130_fd_sc_hd__o211ai_2 _0732_ (.A1(_0269_),
    .A2(_0270_),
    .B1(_0278_),
    .C1(_0279_),
    .Y(_0281_));
 sky130_fd_sc_hd__nand2_1 _0733_ (.A(_0280_),
    .B(_0281_),
    .Y(_0282_));
 sky130_fd_sc_hd__a21oi_1 _0734_ (.A1(_0280_),
    .A2(_0281_),
    .B1(_0126_),
    .Y(_0283_));
 sky130_fd_sc_hd__and3_1 _0735_ (.A(_0126_),
    .B(_0280_),
    .C(_0281_),
    .X(_0284_));
 sky130_fd_sc_hd__a22o_1 _0736_ (.A1(net2),
    .A2(net5),
    .B1(_0088_),
    .B2(_0150_),
    .X(_0285_));
 sky130_fd_sc_hd__a21oi_1 _0737_ (.A1(_0146_),
    .A2(_0189_),
    .B1(_0285_),
    .Y(_0286_));
 sky130_fd_sc_hd__and3_1 _0738_ (.A(_0146_),
    .B(_0189_),
    .C(_0285_),
    .X(_0287_));
 sky130_fd_sc_hd__or2_1 _0739_ (.A(_0286_),
    .B(_0287_),
    .X(_0288_));
 sky130_fd_sc_hd__or3_1 _0740_ (.A(net13),
    .B(_0286_),
    .C(_0287_),
    .X(_0289_));
 sky130_fd_sc_hd__o21bai_2 _0741_ (.A1(_0284_),
    .A2(_0289_),
    .B1_N(_0283_),
    .Y(_0290_));
 sky130_fd_sc_hd__xor2_1 _0742_ (.A(_0170_),
    .B(_0282_),
    .X(_0291_));
 sky130_fd_sc_hd__xnor2_2 _0743_ (.A(_0290_),
    .B(_0291_),
    .Y(_0292_));
 sky130_fd_sc_hd__xnor2_4 _0744_ (.A(_0277_),
    .B(_0292_),
    .Y(_0293_));
 sky130_fd_sc_hd__nand2_1 _0745_ (.A(_0232_),
    .B(_0293_),
    .Y(_0294_));
 sky130_fd_sc_hd__or4_1 _0746_ (.A(net12),
    .B(_0180_),
    .C(_0286_),
    .D(_0287_),
    .X(_0295_));
 sky130_fd_sc_hd__o31ai_2 _0747_ (.A1(net12),
    .A2(_0286_),
    .A3(_0287_),
    .B1(_0180_),
    .Y(_0296_));
 sky130_fd_sc_hd__a211o_1 _0748_ (.A1(_0295_),
    .A2(_0296_),
    .B1(_0283_),
    .C1(_0284_),
    .X(_0297_));
 sky130_fd_sc_hd__o211ai_2 _0749_ (.A1(_0283_),
    .A2(_0284_),
    .B1(_0295_),
    .C1(_0296_),
    .Y(_0298_));
 sky130_fd_sc_hd__nand2_1 _0750_ (.A(_0297_),
    .B(_0298_),
    .Y(_0299_));
 sky130_fd_sc_hd__nand3_1 _0751_ (.A(_0179_),
    .B(_0297_),
    .C(_0298_),
    .Y(_0300_));
 sky130_fd_sc_hd__o21bai_1 _0752_ (.A1(_0267_),
    .A2(_0272_),
    .B1_N(_0266_),
    .Y(_0301_));
 sky130_fd_sc_hd__or2_1 _0753_ (.A(net5),
    .B(net4),
    .X(_0302_));
 sky130_fd_sc_hd__nand2_1 _0754_ (.A(net5),
    .B(net4),
    .Y(_0303_));
 sky130_fd_sc_hd__and3_1 _0755_ (.A(net19),
    .B(_0302_),
    .C(_0303_),
    .X(_0304_));
 sky130_fd_sc_hd__xor2_1 _0756_ (.A(_0162_),
    .B(_0304_),
    .X(_0305_));
 sky130_fd_sc_hd__xnor2_2 _0757_ (.A(_0301_),
    .B(_0305_),
    .Y(_0306_));
 sky130_fd_sc_hd__xnor2_4 _0758_ (.A(_0087_),
    .B(_0306_),
    .Y(_0307_));
 sky130_fd_sc_hd__nand2_1 _0759_ (.A(_0088_),
    .B(_0143_),
    .Y(_0308_));
 sky130_fd_sc_hd__nand2_1 _0760_ (.A(_0271_),
    .B(_0308_),
    .Y(_0309_));
 sky130_fd_sc_hd__xnor2_2 _0761_ (.A(_0288_),
    .B(_0309_),
    .Y(_0310_));
 sky130_fd_sc_hd__xnor2_4 _0762_ (.A(_0307_),
    .B(_0310_),
    .Y(_0311_));
 sky130_fd_sc_hd__a21o_1 _0763_ (.A1(_0297_),
    .A2(_0298_),
    .B1(_0179_),
    .X(_0312_));
 sky130_fd_sc_hd__nand2_1 _0764_ (.A(net13),
    .B(_0312_),
    .Y(_0313_));
 sky130_fd_sc_hd__o21ai_1 _0765_ (.A1(_0311_),
    .A2(_0313_),
    .B1(_0300_),
    .Y(_0314_));
 sky130_fd_sc_hd__or2_1 _0766_ (.A(_0232_),
    .B(_0293_),
    .X(_0315_));
 sky130_fd_sc_hd__xnor2_1 _0767_ (.A(_0232_),
    .B(_0293_),
    .Y(_0316_));
 sky130_fd_sc_hd__a21bo_2 _0768_ (.A1(_0314_),
    .A2(_0315_),
    .B1_N(_0294_),
    .X(_0317_));
 sky130_fd_sc_hd__xor2_1 _0769_ (.A(_0256_),
    .B(_0307_),
    .X(_0318_));
 sky130_fd_sc_hd__xnor2_2 _0770_ (.A(_0293_),
    .B(_0318_),
    .Y(_0319_));
 sky130_fd_sc_hd__mux2_1 _0771_ (.A0(_0163_),
    .A1(_0256_),
    .S(\start_seg[0] ),
    .X(_0320_));
 sky130_fd_sc_hd__xor2_1 _0772_ (.A(_0150_),
    .B(_0320_),
    .X(_0321_));
 sky130_fd_sc_hd__nand3_1 _0773_ (.A(_0110_),
    .B(_0276_),
    .C(_0290_),
    .Y(_0322_));
 sky130_fd_sc_hd__or3_1 _0774_ (.A(_0110_),
    .B(_0276_),
    .C(_0290_),
    .X(_0323_));
 sky130_fd_sc_hd__and2_1 _0775_ (.A(_0322_),
    .B(_0323_),
    .X(_0324_));
 sky130_fd_sc_hd__xnor2_1 _0776_ (.A(_0307_),
    .B(_0321_),
    .Y(_0325_));
 sky130_fd_sc_hd__xnor2_1 _0777_ (.A(_0324_),
    .B(_0325_),
    .Y(_0326_));
 sky130_fd_sc_hd__xor2_2 _0778_ (.A(_0319_),
    .B(_0326_),
    .X(_0327_));
 sky130_fd_sc_hd__xnor2_4 _0779_ (.A(_0317_),
    .B(_0327_),
    .Y(_0328_));
 sky130_fd_sc_hd__xnor2_1 _0780_ (.A(net13),
    .B(_0311_),
    .Y(_0329_));
 sky130_fd_sc_hd__xnor2_1 _0781_ (.A(_0089_),
    .B(_0321_),
    .Y(_0330_));
 sky130_fd_sc_hd__a21oi_1 _0782_ (.A1(_0322_),
    .A2(_0323_),
    .B1(_0330_),
    .Y(_0331_));
 sky130_fd_sc_hd__and3_1 _0783_ (.A(_0322_),
    .B(_0323_),
    .C(_0330_),
    .X(_0332_));
 sky130_fd_sc_hd__or2_1 _0784_ (.A(_0331_),
    .B(_0332_),
    .X(_0333_));
 sky130_fd_sc_hd__or3_1 _0785_ (.A(_0143_),
    .B(_0331_),
    .C(_0332_),
    .X(_0334_));
 sky130_fd_sc_hd__xnor2_1 _0786_ (.A(_0329_),
    .B(_0333_),
    .Y(_0335_));
 sky130_fd_sc_hd__xnor2_1 _0787_ (.A(_0328_),
    .B(_0335_),
    .Y(_0336_));
 sky130_fd_sc_hd__nand2_2 _0788_ (.A(_0143_),
    .B(_0336_),
    .Y(_0337_));
 sky130_fd_sc_hd__or2_1 _0789_ (.A(_0143_),
    .B(_0336_),
    .X(_0338_));
 sky130_fd_sc_hd__and2_1 _0790_ (.A(_0337_),
    .B(_0338_),
    .X(_0339_));
 sky130_fd_sc_hd__xnor2_1 _0791_ (.A(_0220_),
    .B(_0319_),
    .Y(_0340_));
 sky130_fd_sc_hd__xnor2_2 _0792_ (.A(_0317_),
    .B(_0340_),
    .Y(_0341_));
 sky130_fd_sc_hd__a21o_1 _0793_ (.A1(_0300_),
    .A2(_0312_),
    .B1(_0282_),
    .X(_0342_));
 sky130_fd_sc_hd__nand3_1 _0794_ (.A(_0282_),
    .B(_0300_),
    .C(_0312_),
    .Y(_0343_));
 sky130_fd_sc_hd__o211ai_1 _0795_ (.A1(net14),
    .A2(_0311_),
    .B1(_0342_),
    .C1(_0343_),
    .Y(_0344_));
 sky130_fd_sc_hd__a211o_1 _0796_ (.A1(_0342_),
    .A2(_0343_),
    .B1(net13),
    .C1(_0311_),
    .X(_0345_));
 sky130_fd_sc_hd__a2bb2oi_1 _0797_ (.A1_N(net13),
    .A2_N(_0311_),
    .B1(_0342_),
    .B2(_0343_),
    .Y(_0346_));
 sky130_fd_sc_hd__and4bb_1 _0798_ (.A_N(net13),
    .B_N(_0311_),
    .C(_0342_),
    .D(_0343_),
    .X(_0347_));
 sky130_fd_sc_hd__or2_1 _0799_ (.A(_0346_),
    .B(_0347_),
    .X(_0348_));
 sky130_fd_sc_hd__or3_1 _0800_ (.A(net15),
    .B(_0346_),
    .C(_0347_),
    .X(_0349_));
 sky130_fd_sc_hd__o21ai_1 _0801_ (.A1(_0346_),
    .A2(_0347_),
    .B1(net15),
    .Y(_0350_));
 sky130_fd_sc_hd__a311o_1 _0802_ (.A1(net15),
    .A2(_0344_),
    .A3(_0345_),
    .B1(net13),
    .C1(_0333_),
    .X(_0351_));
 sky130_fd_sc_hd__a21oi_1 _0803_ (.A1(_0349_),
    .A2(_0351_),
    .B1(_0200_),
    .Y(_0352_));
 sky130_fd_sc_hd__xnor2_1 _0804_ (.A(_0314_),
    .B(_0316_),
    .Y(_0353_));
 sky130_fd_sc_hd__xnor2_1 _0805_ (.A(_0275_),
    .B(_0299_),
    .Y(_0354_));
 sky130_fd_sc_hd__xnor2_2 _0806_ (.A(_0353_),
    .B(_0354_),
    .Y(_0355_));
 sky130_fd_sc_hd__and3_1 _0807_ (.A(_0200_),
    .B(_0349_),
    .C(_0351_),
    .X(_0356_));
 sky130_fd_sc_hd__mux2_2 _0808_ (.A0(_0356_),
    .A1(_0352_),
    .S(_0355_),
    .X(_0357_));
 sky130_fd_sc_hd__xnor2_4 _0809_ (.A(_0341_),
    .B(_0357_),
    .Y(_0358_));
 sky130_fd_sc_hd__xor2_4 _0810_ (.A(_0328_),
    .B(_0358_),
    .X(_0359_));
 sky130_fd_sc_hd__xor2_4 _0811_ (.A(_0311_),
    .B(_0359_),
    .X(_0360_));
 sky130_fd_sc_hd__xnor2_1 _0812_ (.A(_0339_),
    .B(_0360_),
    .Y(_0361_));
 sky130_fd_sc_hd__xor2_1 _0813_ (.A(_0293_),
    .B(_0348_),
    .X(_0362_));
 sky130_fd_sc_hd__xnor2_1 _0814_ (.A(_0355_),
    .B(_0362_),
    .Y(_0363_));
 sky130_fd_sc_hd__nor2_1 _0815_ (.A(_0352_),
    .B(_0356_),
    .Y(_0364_));
 sky130_fd_sc_hd__xnor2_2 _0816_ (.A(_0363_),
    .B(_0364_),
    .Y(_0365_));
 sky130_fd_sc_hd__xor2_1 _0817_ (.A(_0299_),
    .B(_0334_),
    .X(_0366_));
 sky130_fd_sc_hd__a21oi_1 _0818_ (.A1(_0349_),
    .A2(_0350_),
    .B1(_0366_),
    .Y(_0367_));
 sky130_fd_sc_hd__and3_1 _0819_ (.A(_0349_),
    .B(_0350_),
    .C(_0366_),
    .X(_0368_));
 sky130_fd_sc_hd__nor2_2 _0820_ (.A(_0367_),
    .B(_0368_),
    .Y(_0369_));
 sky130_fd_sc_hd__o211a_1 _0821_ (.A1(_0178_),
    .A2(_0369_),
    .B1(_0336_),
    .C1(net13),
    .X(_0370_));
 sky130_fd_sc_hd__a21oi_1 _0822_ (.A1(_0178_),
    .A2(_0369_),
    .B1(_0370_),
    .Y(_0371_));
 sky130_fd_sc_hd__mux2_1 _0823_ (.A0(_0365_),
    .A1(_0105_),
    .S(_0371_),
    .X(_0372_));
 sky130_fd_sc_hd__o21ba_1 _0824_ (.A1(_0105_),
    .A2(_0365_),
    .B1_N(_0372_),
    .X(_0373_));
 sky130_fd_sc_hd__xor2_1 _0825_ (.A(_0196_),
    .B(_0359_),
    .X(_0374_));
 sky130_fd_sc_hd__xnor2_1 _0826_ (.A(_0373_),
    .B(_0374_),
    .Y(_0375_));
 sky130_fd_sc_hd__or3_1 _0827_ (.A(mode_dec),
    .B(_0361_),
    .C(_0375_),
    .X(_0376_));
 sky130_fd_sc_hd__a21oi_1 _0828_ (.A1(_0083_),
    .A2(_0375_),
    .B1(_0086_),
    .Y(_0377_));
 sky130_fd_sc_hd__o21bai_1 _0829_ (.A1(_0086_),
    .A2(_0361_),
    .B1_N(_0377_),
    .Y(_0378_));
 sky130_fd_sc_hd__o211a_2 _0830_ (.A1(_0083_),
    .A2(_0265_),
    .B1(_0376_),
    .C1(_0378_),
    .X(uo_out[0]));
 sky130_fd_sc_hd__xnor2_1 _0831_ (.A(_0179_),
    .B(_0369_),
    .Y(_0379_));
 sky130_fd_sc_hd__xnor2_2 _0832_ (.A(_0348_),
    .B(_0379_),
    .Y(_0380_));
 sky130_fd_sc_hd__xnor2_4 _0833_ (.A(_0337_),
    .B(_0380_),
    .Y(_0381_));
 sky130_fd_sc_hd__or2_1 _0834_ (.A(net15),
    .B(_0381_),
    .X(_0382_));
 sky130_fd_sc_hd__nand2_1 _0835_ (.A(_0125_),
    .B(_0381_),
    .Y(_0383_));
 sky130_fd_sc_hd__and2_1 _0836_ (.A(_0382_),
    .B(_0383_),
    .X(_0384_));
 sky130_fd_sc_hd__xnor2_1 _0837_ (.A(_0369_),
    .B(_0384_),
    .Y(_0385_));
 sky130_fd_sc_hd__a21oi_1 _0838_ (.A1(net13),
    .A2(_0360_),
    .B1(_0385_),
    .Y(_0386_));
 sky130_fd_sc_hd__a31o_1 _0839_ (.A1(net13),
    .A2(_0360_),
    .A3(_0385_),
    .B1(mode_dec),
    .X(_0387_));
 sky130_fd_sc_hd__nor2_1 _0840_ (.A(net14),
    .B(_0168_),
    .Y(_0388_));
 sky130_fd_sc_hd__or2_1 _0841_ (.A(_0233_),
    .B(_0388_),
    .X(_0389_));
 sky130_fd_sc_hd__nor2_1 _0842_ (.A(net14),
    .B(_0244_),
    .Y(_0390_));
 sky130_fd_sc_hd__inv_2 _0843_ (.A(_0390_),
    .Y(_0391_));
 sky130_fd_sc_hd__xnor2_1 _0844_ (.A(_0244_),
    .B(_0389_),
    .Y(_0392_));
 sky130_fd_sc_hd__or3_1 _0845_ (.A(_0228_),
    .B(_0229_),
    .C(_0392_),
    .X(_0393_));
 sky130_fd_sc_hd__o21ai_1 _0846_ (.A1(_0228_),
    .A2(_0229_),
    .B1(_0392_),
    .Y(_0394_));
 sky130_fd_sc_hd__a21oi_1 _0847_ (.A1(_0241_),
    .A2(_0242_),
    .B1(_0211_),
    .Y(_0395_));
 sky130_fd_sc_hd__and3_1 _0848_ (.A(_0211_),
    .B(_0241_),
    .C(_0242_),
    .X(_0396_));
 sky130_fd_sc_hd__or3_1 _0849_ (.A(_0391_),
    .B(_0395_),
    .C(_0396_),
    .X(_0397_));
 sky130_fd_sc_hd__o21ai_1 _0850_ (.A1(_0395_),
    .A2(_0396_),
    .B1(_0391_),
    .Y(_0398_));
 sky130_fd_sc_hd__nand2_1 _0851_ (.A(_0397_),
    .B(_0398_),
    .Y(_0399_));
 sky130_fd_sc_hd__and3_1 _0852_ (.A(net15),
    .B(_0397_),
    .C(_0398_),
    .X(_0400_));
 sky130_fd_sc_hd__nand3_1 _0853_ (.A(net15),
    .B(_0397_),
    .C(_0398_),
    .Y(_0401_));
 sky130_fd_sc_hd__a21o_1 _0854_ (.A1(_0397_),
    .A2(_0398_),
    .B1(net15),
    .X(_0402_));
 sky130_fd_sc_hd__and4_1 _0855_ (.A(net14),
    .B(_0239_),
    .C(_0393_),
    .D(_0394_),
    .X(_0403_));
 sky130_fd_sc_hd__a31oi_1 _0856_ (.A1(net14),
    .A2(_0393_),
    .A3(_0394_),
    .B1(_0239_),
    .Y(_0404_));
 sky130_fd_sc_hd__a211o_1 _0857_ (.A1(_0401_),
    .A2(_0402_),
    .B1(_0403_),
    .C1(_0404_),
    .X(_0405_));
 sky130_fd_sc_hd__o211ai_1 _0858_ (.A1(_0403_),
    .A2(_0404_),
    .B1(_0401_),
    .C1(_0402_),
    .Y(_0406_));
 sky130_fd_sc_hd__and2_1 _0859_ (.A(_0405_),
    .B(_0406_),
    .X(_0407_));
 sky130_fd_sc_hd__or2_1 _0860_ (.A(_0083_),
    .B(_0407_),
    .X(_0408_));
 sky130_fd_sc_hd__o211a_4 _0861_ (.A1(_0386_),
    .A2(_0387_),
    .B1(_0408_),
    .C1(net19),
    .X(uo_out[1]));
 sky130_fd_sc_hd__xnor2_1 _0862_ (.A(_0106_),
    .B(_0365_),
    .Y(_0409_));
 sky130_fd_sc_hd__xnor2_1 _0863_ (.A(_0355_),
    .B(_0369_),
    .Y(_0410_));
 sky130_fd_sc_hd__xnor2_1 _0864_ (.A(_0371_),
    .B(_0410_),
    .Y(_0411_));
 sky130_fd_sc_hd__xnor2_2 _0865_ (.A(_0409_),
    .B(_0411_),
    .Y(_0412_));
 sky130_fd_sc_hd__nor2_1 _0866_ (.A(_0110_),
    .B(_0412_),
    .Y(_0413_));
 sky130_fd_sc_hd__xor2_1 _0867_ (.A(_0110_),
    .B(_0412_),
    .X(_0414_));
 sky130_fd_sc_hd__a22o_1 _0868_ (.A1(net12),
    .A2(_0360_),
    .B1(_0381_),
    .B2(net15),
    .X(_0415_));
 sky130_fd_sc_hd__nand2_1 _0869_ (.A(_0382_),
    .B(_0415_),
    .Y(_0416_));
 sky130_fd_sc_hd__xnor2_1 _0870_ (.A(_0414_),
    .B(_0416_),
    .Y(_0417_));
 sky130_fd_sc_hd__xnor2_1 _0871_ (.A(_0365_),
    .B(_0381_),
    .Y(_0418_));
 sky130_fd_sc_hd__nand2_1 _0872_ (.A(_0417_),
    .B(_0418_),
    .Y(_0419_));
 sky130_fd_sc_hd__o21a_1 _0873_ (.A1(_0417_),
    .A2(_0418_),
    .B1(_0083_),
    .X(_0420_));
 sky130_fd_sc_hd__nand2b_1 _0874_ (.A_N(_0246_),
    .B(_0252_),
    .Y(_0421_));
 sky130_fd_sc_hd__xnor2_1 _0875_ (.A(_0205_),
    .B(_0238_),
    .Y(_0422_));
 sky130_fd_sc_hd__a21o_1 _0876_ (.A1(_0249_),
    .A2(_0250_),
    .B1(_0422_),
    .X(_0423_));
 sky130_fd_sc_hd__nand3_1 _0877_ (.A(_0249_),
    .B(_0250_),
    .C(_0422_),
    .Y(_0424_));
 sky130_fd_sc_hd__nand3_2 _0878_ (.A(_0421_),
    .B(_0423_),
    .C(_0424_),
    .Y(_0425_));
 sky130_fd_sc_hd__a21o_1 _0879_ (.A1(_0423_),
    .A2(_0424_),
    .B1(_0421_),
    .X(_0426_));
 sky130_fd_sc_hd__nand2_1 _0880_ (.A(_0425_),
    .B(_0426_),
    .Y(_0427_));
 sky130_fd_sc_hd__nand3b_1 _0881_ (.A_N(_0110_),
    .B(_0425_),
    .C(_0426_),
    .Y(_0428_));
 sky130_fd_sc_hd__a21bo_1 _0882_ (.A1(_0425_),
    .A2(_0426_),
    .B1_N(_0110_),
    .X(_0429_));
 sky130_fd_sc_hd__a41o_1 _0883_ (.A1(net12),
    .A2(_0393_),
    .A3(_0394_),
    .A4(_0402_),
    .B1(_0400_),
    .X(_0430_));
 sky130_fd_sc_hd__nand3_1 _0884_ (.A(_0428_),
    .B(_0429_),
    .C(_0430_),
    .Y(_0431_));
 sky130_fd_sc_hd__a21o_1 _0885_ (.A1(_0428_),
    .A2(_0429_),
    .B1(_0430_),
    .X(_0432_));
 sky130_fd_sc_hd__xor2_1 _0886_ (.A(_0251_),
    .B(_0399_),
    .X(_0433_));
 sky130_fd_sc_hd__a21boi_1 _0887_ (.A1(_0431_),
    .A2(_0432_),
    .B1_N(_0433_),
    .Y(_0434_));
 sky130_fd_sc_hd__and3b_1 _0888_ (.A_N(_0433_),
    .B(_0432_),
    .C(_0431_),
    .X(_0435_));
 sky130_fd_sc_hd__nor2_1 _0889_ (.A(_0434_),
    .B(_0435_),
    .Y(_0436_));
 sky130_fd_sc_hd__a221oi_4 _0890_ (.A1(_0419_),
    .A2(_0420_),
    .B1(_0436_),
    .B2(mode_dec),
    .C1(_0086_),
    .Y(uo_out[2]));
 sky130_fd_sc_hd__a31o_1 _0891_ (.A1(_0382_),
    .A2(_0414_),
    .A3(_0415_),
    .B1(_0413_),
    .X(_0437_));
 sky130_fd_sc_hd__xor2_1 _0892_ (.A(_0165_),
    .B(_0358_),
    .X(_0438_));
 sky130_fd_sc_hd__xnor2_1 _0893_ (.A(_0412_),
    .B(_0438_),
    .Y(_0439_));
 sky130_fd_sc_hd__xnor2_1 _0894_ (.A(_0375_),
    .B(_0439_),
    .Y(_0440_));
 sky130_fd_sc_hd__nor2_1 _0895_ (.A(_0437_),
    .B(_0440_),
    .Y(_0441_));
 sky130_fd_sc_hd__a21o_1 _0896_ (.A1(_0437_),
    .A2(_0440_),
    .B1(mode_dec),
    .X(_0442_));
 sky130_fd_sc_hd__a21bo_1 _0897_ (.A1(_0428_),
    .A2(_0430_),
    .B1_N(_0429_),
    .X(_0443_));
 sky130_fd_sc_hd__a21oi_1 _0898_ (.A1(_0425_),
    .A2(_0426_),
    .B1(_0320_),
    .Y(_0444_));
 sky130_fd_sc_hd__and3_1 _0899_ (.A(_0320_),
    .B(_0425_),
    .C(_0426_),
    .X(_0445_));
 sky130_fd_sc_hd__o211a_1 _0900_ (.A1(_0444_),
    .A2(_0445_),
    .B1(_0261_),
    .C1(_0262_),
    .X(_0446_));
 sky130_fd_sc_hd__a211oi_1 _0901_ (.A1(_0261_),
    .A2(_0262_),
    .B1(_0444_),
    .C1(_0445_),
    .Y(_0447_));
 sky130_fd_sc_hd__or3_1 _0902_ (.A(_0443_),
    .B(_0446_),
    .C(_0447_),
    .X(_0448_));
 sky130_fd_sc_hd__o21ai_1 _0903_ (.A1(_0446_),
    .A2(_0447_),
    .B1(_0443_),
    .Y(_0449_));
 sky130_fd_sc_hd__nand2_1 _0904_ (.A(_0448_),
    .B(_0449_),
    .Y(_0450_));
 sky130_fd_sc_hd__nand2_1 _0905_ (.A(mode_dec),
    .B(_0450_),
    .Y(_0451_));
 sky130_fd_sc_hd__o211a_4 _0906_ (.A1(_0441_),
    .A2(_0442_),
    .B1(_0451_),
    .C1(net19),
    .X(uo_out[3]));
 sky130_fd_sc_hd__xnor2_1 _0907_ (.A(_0244_),
    .B(_0260_),
    .Y(_0452_));
 sky130_fd_sc_hd__nor2_1 _0908_ (.A(_0450_),
    .B(_0452_),
    .Y(_0453_));
 sky130_fd_sc_hd__a21o_1 _0909_ (.A1(_0450_),
    .A2(_0452_),
    .B1(_0083_),
    .X(_0454_));
 sky130_fd_sc_hd__o221a_4 _0910_ (.A1(mode_dec),
    .A2(_0360_),
    .B1(_0453_),
    .B2(_0454_),
    .C1(net19),
    .X(uo_out[4]));
 sky130_fd_sc_hd__and3_1 _0911_ (.A(net12),
    .B(_0263_),
    .C(_0264_),
    .X(_0455_));
 sky130_fd_sc_hd__a21o_1 _0912_ (.A1(_0405_),
    .A2(_0406_),
    .B1(_0178_),
    .X(_0456_));
 sky130_fd_sc_hd__and3_1 _0913_ (.A(_0178_),
    .B(_0405_),
    .C(_0406_),
    .X(_0457_));
 sky130_fd_sc_hd__nand2_1 _0914_ (.A(_0178_),
    .B(_0407_),
    .Y(_0458_));
 sky130_fd_sc_hd__a21oi_1 _0915_ (.A1(_0456_),
    .A2(_0458_),
    .B1(_0399_),
    .Y(_0459_));
 sky130_fd_sc_hd__and3_1 _0916_ (.A(_0399_),
    .B(_0456_),
    .C(_0458_),
    .X(_0460_));
 sky130_fd_sc_hd__nor2_1 _0917_ (.A(_0459_),
    .B(_0460_),
    .Y(_0461_));
 sky130_fd_sc_hd__nor2_1 _0918_ (.A(_0455_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__a21o_1 _0919_ (.A1(_0455_),
    .A2(_0461_),
    .B1(_0083_),
    .X(_0463_));
 sky130_fd_sc_hd__o221a_4 _0920_ (.A1(mode_dec),
    .A2(_0381_),
    .B1(_0462_),
    .B2(_0463_),
    .C1(net19),
    .X(uo_out[5]));
 sky130_fd_sc_hd__xnor2_1 _0921_ (.A(_0407_),
    .B(_0427_),
    .Y(_0464_));
 sky130_fd_sc_hd__a41oi_2 _0922_ (.A1(net14),
    .A2(_0263_),
    .A3(_0264_),
    .A4(_0456_),
    .B1(_0457_),
    .Y(_0465_));
 sky130_fd_sc_hd__xnor2_1 _0923_ (.A(_0106_),
    .B(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__xnor2_1 _0924_ (.A(_0436_),
    .B(_0466_),
    .Y(_0467_));
 sky130_fd_sc_hd__nor2_1 _0925_ (.A(_0464_),
    .B(_0467_),
    .Y(_0468_));
 sky130_fd_sc_hd__a21o_1 _0926_ (.A1(_0464_),
    .A2(_0467_),
    .B1(_0083_),
    .X(_0469_));
 sky130_fd_sc_hd__a21oi_1 _0927_ (.A1(_0083_),
    .A2(_0412_),
    .B1(_0086_),
    .Y(_0470_));
 sky130_fd_sc_hd__o21a_2 _0928_ (.A1(_0468_),
    .A2(_0469_),
    .B1(_0470_),
    .X(uo_out[6]));
 sky130_fd_sc_hd__xnor2_1 _0929_ (.A(_0162_),
    .B(_0260_),
    .Y(_0471_));
 sky130_fd_sc_hd__xnor2_1 _0930_ (.A(_0450_),
    .B(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__o211ai_1 _0931_ (.A1(_0434_),
    .A2(_0435_),
    .B1(_0465_),
    .C1(_0105_),
    .Y(_0473_));
 sky130_fd_sc_hd__or4_1 _0932_ (.A(_0105_),
    .B(_0434_),
    .C(_0435_),
    .D(_0465_),
    .X(_0474_));
 sky130_fd_sc_hd__nand2_1 _0933_ (.A(_0473_),
    .B(_0474_),
    .Y(_0475_));
 sky130_fd_sc_hd__xnor2_1 _0934_ (.A(_0472_),
    .B(_0475_),
    .Y(_0476_));
 sky130_fd_sc_hd__o21a_4 _0935_ (.A1(_0083_),
    .A2(_0476_),
    .B1(_0377_),
    .X(uo_out[7]));
 sky130_fd_sc_hd__and2b_1 _0936_ (.A_N(net20),
    .B(\sys_state[0] ),
    .X(_0477_));
 sky130_fd_sc_hd__nand2b_1 _0937_ (.A_N(net20),
    .B(\sys_state[0] ),
    .Y(_0478_));
 sky130_fd_sc_hd__nor2_1 _0938_ (.A(net127),
    .B(_0478_),
    .Y(_0000_));
 sky130_fd_sc_hd__and2_1 _0939_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .X(_0479_));
 sky130_fd_sc_hd__nand2_1 _0940_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .Y(_0480_));
 sky130_fd_sc_hd__nor2_1 _0941_ (.A(\counter[0] ),
    .B(\counter[1] ),
    .Y(_0481_));
 sky130_fd_sc_hd__and3b_1 _0942_ (.A_N(_0481_),
    .B(_0477_),
    .C(_0480_),
    .X(_0001_));
 sky130_fd_sc_hd__or2_1 _0943_ (.A(net22),
    .B(_0479_),
    .X(_0482_));
 sky130_fd_sc_hd__nand2_1 _0944_ (.A(net22),
    .B(_0479_),
    .Y(_0483_));
 sky130_fd_sc_hd__and3_1 _0945_ (.A(_0477_),
    .B(_0482_),
    .C(_0483_),
    .X(_0002_));
 sky130_fd_sc_hd__a31o_1 _0946_ (.A1(\counter[0] ),
    .A2(\counter[1] ),
    .A3(net22),
    .B1(\counter[3] ),
    .X(_0484_));
 sky130_fd_sc_hd__nor2_1 _0947_ (.A(\counter[3] ),
    .B(_0478_),
    .Y(_0485_));
 sky130_fd_sc_hd__or2_2 _0948_ (.A(\counter[3] ),
    .B(_0478_),
    .X(_0486_));
 sky130_fd_sc_hd__nand3_1 _0949_ (.A(net22),
    .B(\counter[3] ),
    .C(_0479_),
    .Y(_0487_));
 sky130_fd_sc_hd__and3_1 _0950_ (.A(_0477_),
    .B(_0484_),
    .C(_0487_),
    .X(_0003_));
 sky130_fd_sc_hd__and2_1 _0951_ (.A(\counter[3] ),
    .B(_0477_),
    .X(_0488_));
 sky130_fd_sc_hd__nand2_2 _0952_ (.A(\counter[3] ),
    .B(_0477_),
    .Y(_0489_));
 sky130_fd_sc_hd__nand2b_1 _0953_ (.A_N(net21),
    .B(\counter[2] ),
    .Y(_0490_));
 sky130_fd_sc_hd__or3_4 _0954_ (.A(net21),
    .B(_0483_),
    .C(_0489_),
    .X(_0491_));
 sky130_fd_sc_hd__inv_2 _0955_ (.A(_0491_),
    .Y(_0492_));
 sky130_fd_sc_hd__a31o_1 _0956_ (.A1(net21),
    .A2(_0477_),
    .A3(_0487_),
    .B1(_0492_),
    .X(_0004_));
 sky130_fd_sc_hd__or4_1 _0957_ (.A(net35),
    .B(net29),
    .C(net8),
    .D(net33),
    .X(_0493_));
 sky130_fd_sc_hd__nor3_1 _0958_ (.A(net20),
    .B(\sys_state[0] ),
    .C(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__nand2_1 _0959_ (.A(net2),
    .B(net3),
    .Y(_0495_));
 sky130_fd_sc_hd__a21oi_1 _0960_ (.A1(_0078_),
    .A2(_0081_),
    .B1(_0302_),
    .Y(_0496_));
 sky130_fd_sc_hd__and3_1 _0961_ (.A(_0494_),
    .B(_0495_),
    .C(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__or2_1 _0962_ (.A(net21),
    .B(_0487_),
    .X(_0498_));
 sky130_fd_sc_hd__a221o_1 _0963_ (.A1(_0084_),
    .A2(net18),
    .B1(_0477_),
    .B2(_0498_),
    .C1(_0497_),
    .X(\sys_next_state[0] ));
 sky130_fd_sc_hd__nor2_1 _0964_ (.A(net2),
    .B(_0302_),
    .Y(_0499_));
 sky130_fd_sc_hd__a2bb2o_1 _0965_ (.A1_N(_0303_),
    .A2_N(_0495_),
    .B1(_0499_),
    .B2(net3),
    .X(_0500_));
 sky130_fd_sc_hd__a22o_1 _0966_ (.A1(_0084_),
    .A2(net18),
    .B1(_0494_),
    .B2(_0500_),
    .X(\sys_next_state[1] ));
 sky130_fd_sc_hd__nand2b_4 _0967_ (.A_N(\sys_state[0] ),
    .B(\sys_state[1] ),
    .Y(_0501_));
 sky130_fd_sc_hd__mux2_1 _0968_ (.A0(net2),
    .A1(\start_seg[0] ),
    .S(_0501_),
    .X(_0005_));
 sky130_fd_sc_hd__mux2_1 _0969_ (.A0(net3),
    .A1(\start_seg[1] ),
    .S(_0501_),
    .X(_0006_));
 sky130_fd_sc_hd__and3b_1 _0970_ (.A_N(\sys_state[0] ),
    .B(net4),
    .C(net20),
    .X(_0502_));
 sky130_fd_sc_hd__a21o_1 _0971_ (.A1(\start_seg[2] ),
    .A2(_0501_),
    .B1(_0502_),
    .X(_0007_));
 sky130_fd_sc_hd__mux2_1 _0972_ (.A0(net5),
    .A1(\start_seg[3] ),
    .S(_0501_),
    .X(_0008_));
 sky130_fd_sc_hd__mux2_1 _0973_ (.A0(mode_dec),
    .A1(net10),
    .S(_0086_),
    .X(_0009_));
 sky130_fd_sc_hd__mux2_1 _0974_ (.A0(_0086_),
    .A1(net20),
    .S(net27),
    .X(_0503_));
 sky130_fd_sc_hd__o21ai_1 _0975_ (.A1(_0078_),
    .A2(_0501_),
    .B1(_0503_),
    .Y(_0010_));
 sky130_fd_sc_hd__a21oi_1 _0976_ (.A1(\sys_state[1] ),
    .A2(net27),
    .B1(net25),
    .Y(_0504_));
 sky130_fd_sc_hd__and3_1 _0977_ (.A(\sys_state[1] ),
    .B(net27),
    .C(net25),
    .X(_0505_));
 sky130_fd_sc_hd__nor2_1 _0978_ (.A(_0504_),
    .B(_0505_),
    .Y(_0506_));
 sky130_fd_sc_hd__mux2_1 _0979_ (.A0(net3),
    .A1(_0506_),
    .S(_0501_),
    .X(_0011_));
 sky130_fd_sc_hd__or2_1 _0980_ (.A(net23),
    .B(_0505_),
    .X(_0507_));
 sky130_fd_sc_hd__nand2_1 _0981_ (.A(net23),
    .B(_0505_),
    .Y(_0508_));
 sky130_fd_sc_hd__a31o_1 _0982_ (.A1(_0501_),
    .A2(_0507_),
    .A3(_0508_),
    .B1(_0502_),
    .X(_0012_));
 sky130_fd_sc_hd__xnor2_1 _0983_ (.A(\curr_seg[3] ),
    .B(_0508_),
    .Y(_0509_));
 sky130_fd_sc_hd__mux2_1 _0984_ (.A0(net5),
    .A1(_0509_),
    .S(_0501_),
    .X(_0013_));
 sky130_fd_sc_hd__mux2_1 _0985_ (.A0(net34),
    .A1(net102),
    .S(_0491_),
    .X(_0014_));
 sky130_fd_sc_hd__mux2_1 _0986_ (.A0(net32),
    .A1(net92),
    .S(_0491_),
    .X(_0015_));
 sky130_fd_sc_hd__mux2_1 _0987_ (.A0(net30),
    .A1(net89),
    .S(_0491_),
    .X(_0016_));
 sky130_fd_sc_hd__mux2_1 _0988_ (.A0(net28),
    .A1(net122),
    .S(_0491_),
    .X(_0017_));
 sky130_fd_sc_hd__or4bb_1 _0989_ (.A(\counter[0] ),
    .B(net21),
    .C_N(net22),
    .D_N(\counter[1] ),
    .X(_0510_));
 sky130_fd_sc_hd__or2_2 _0990_ (.A(_0489_),
    .B(_0510_),
    .X(_0511_));
 sky130_fd_sc_hd__mux2_1 _0991_ (.A0(net34),
    .A1(net114),
    .S(_0511_),
    .X(_0018_));
 sky130_fd_sc_hd__mux2_1 _0992_ (.A0(net32),
    .A1(net121),
    .S(_0511_),
    .X(_0019_));
 sky130_fd_sc_hd__mux2_1 _0993_ (.A0(net30),
    .A1(net100),
    .S(_0511_),
    .X(_0020_));
 sky130_fd_sc_hd__mux2_1 _0994_ (.A0(net28),
    .A1(net90),
    .S(_0511_),
    .X(_0021_));
 sky130_fd_sc_hd__or4b_4 _0995_ (.A(\counter[1] ),
    .B(_0489_),
    .C(_0490_),
    .D_N(\counter[0] ),
    .X(_0512_));
 sky130_fd_sc_hd__mux2_1 _0996_ (.A0(net34),
    .A1(net123),
    .S(_0512_),
    .X(_0022_));
 sky130_fd_sc_hd__mux2_1 _0997_ (.A0(net32),
    .A1(net120),
    .S(_0512_),
    .X(_0023_));
 sky130_fd_sc_hd__mux2_1 _0998_ (.A0(net30),
    .A1(net91),
    .S(_0512_),
    .X(_0024_));
 sky130_fd_sc_hd__mux2_1 _0999_ (.A0(net28),
    .A1(net105),
    .S(_0512_),
    .X(_0025_));
 sky130_fd_sc_hd__and4b_2 _1000_ (.A_N(net21),
    .B(_0481_),
    .C(_0488_),
    .D(net22),
    .X(_0513_));
 sky130_fd_sc_hd__mux2_1 _1001_ (.A0(net88),
    .A1(net34),
    .S(_0513_),
    .X(_0026_));
 sky130_fd_sc_hd__mux2_1 _1002_ (.A0(net82),
    .A1(net32),
    .S(_0513_),
    .X(_0027_));
 sky130_fd_sc_hd__mux2_1 _1003_ (.A0(net83),
    .A1(net30),
    .S(_0513_),
    .X(_0028_));
 sky130_fd_sc_hd__mux2_1 _1004_ (.A0(net110),
    .A1(net28),
    .S(_0513_),
    .X(_0029_));
 sky130_fd_sc_hd__nor2_1 _1005_ (.A(net22),
    .B(net21),
    .Y(_0514_));
 sky130_fd_sc_hd__or3b_2 _1006_ (.A(_0480_),
    .B(_0489_),
    .C_N(_0514_),
    .X(_0515_));
 sky130_fd_sc_hd__mux2_1 _1007_ (.A0(net35),
    .A1(net124),
    .S(_0515_),
    .X(_0030_));
 sky130_fd_sc_hd__mux2_1 _1008_ (.A0(net33),
    .A1(net109),
    .S(_0515_),
    .X(_0031_));
 sky130_fd_sc_hd__mux2_1 _1009_ (.A0(net31),
    .A1(net125),
    .S(_0515_),
    .X(_0032_));
 sky130_fd_sc_hd__mux2_1 _1010_ (.A0(net29),
    .A1(net119),
    .S(_0515_),
    .X(_0033_));
 sky130_fd_sc_hd__or4b_2 _1011_ (.A(\counter[0] ),
    .B(net22),
    .C(net21),
    .D_N(\counter[1] ),
    .X(_0516_));
 sky130_fd_sc_hd__nor2_2 _1012_ (.A(_0489_),
    .B(_0516_),
    .Y(_0517_));
 sky130_fd_sc_hd__mux2_1 _1013_ (.A0(net126),
    .A1(net35),
    .S(_0517_),
    .X(_0034_));
 sky130_fd_sc_hd__mux2_1 _1014_ (.A0(net111),
    .A1(net33),
    .S(_0517_),
    .X(_0035_));
 sky130_fd_sc_hd__mux2_1 _1015_ (.A0(net76),
    .A1(net31),
    .S(_0517_),
    .X(_0036_));
 sky130_fd_sc_hd__mux2_1 _1016_ (.A0(net116),
    .A1(net29),
    .S(_0517_),
    .X(_0037_));
 sky130_fd_sc_hd__or4b_2 _1017_ (.A(\counter[1] ),
    .B(net22),
    .C(net21),
    .D_N(\counter[0] ),
    .X(_0518_));
 sky130_fd_sc_hd__nor2_2 _1018_ (.A(_0489_),
    .B(_0518_),
    .Y(_0519_));
 sky130_fd_sc_hd__mux2_1 _1019_ (.A0(net67),
    .A1(net35),
    .S(_0519_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _1020_ (.A0(net64),
    .A1(net33),
    .S(_0519_),
    .X(_0039_));
 sky130_fd_sc_hd__mux2_1 _1021_ (.A0(net69),
    .A1(net31),
    .S(_0519_),
    .X(_0040_));
 sky130_fd_sc_hd__mux2_1 _1022_ (.A0(net63),
    .A1(net29),
    .S(_0519_),
    .X(_0041_));
 sky130_fd_sc_hd__and3_2 _1023_ (.A(_0481_),
    .B(_0488_),
    .C(_0514_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_1 _1024_ (.A0(net80),
    .A1(net35),
    .S(_0520_),
    .X(_0042_));
 sky130_fd_sc_hd__mux2_1 _1025_ (.A0(net86),
    .A1(net33),
    .S(_0520_),
    .X(_0043_));
 sky130_fd_sc_hd__mux2_1 _1026_ (.A0(net81),
    .A1(net31),
    .S(_0520_),
    .X(_0044_));
 sky130_fd_sc_hd__mux2_1 _1027_ (.A0(net72),
    .A1(net29),
    .S(_0520_),
    .X(_0045_));
 sky130_fd_sc_hd__or3_2 _1028_ (.A(\counter[4] ),
    .B(_0483_),
    .C(_0486_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_1 _1029_ (.A0(net34),
    .A1(net113),
    .S(_0521_),
    .X(_0046_));
 sky130_fd_sc_hd__mux2_1 _1030_ (.A0(net32),
    .A1(net108),
    .S(_0521_),
    .X(_0047_));
 sky130_fd_sc_hd__mux2_1 _1031_ (.A0(net30),
    .A1(net97),
    .S(_0521_),
    .X(_0048_));
 sky130_fd_sc_hd__mux2_1 _1032_ (.A0(net28),
    .A1(net96),
    .S(_0521_),
    .X(_0049_));
 sky130_fd_sc_hd__nor2_2 _1033_ (.A(_0486_),
    .B(_0510_),
    .Y(_0522_));
 sky130_fd_sc_hd__mux2_1 _1034_ (.A0(net107),
    .A1(net34),
    .S(_0522_),
    .X(_0050_));
 sky130_fd_sc_hd__mux2_1 _1035_ (.A0(net112),
    .A1(net32),
    .S(_0522_),
    .X(_0051_));
 sky130_fd_sc_hd__mux2_1 _1036_ (.A0(net66),
    .A1(net30),
    .S(_0522_),
    .X(_0052_));
 sky130_fd_sc_hd__mux2_1 _1037_ (.A0(net68),
    .A1(net28),
    .S(_0522_),
    .X(_0053_));
 sky130_fd_sc_hd__nor4b_1 _1038_ (.A(\counter[1] ),
    .B(_0486_),
    .C(_0490_),
    .D_N(\counter[0] ),
    .Y(_0523_));
 sky130_fd_sc_hd__mux2_1 _1039_ (.A0(net70),
    .A1(net34),
    .S(net17),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _1040_ (.A0(net93),
    .A1(net32),
    .S(net17),
    .X(_0055_));
 sky130_fd_sc_hd__mux2_1 _1041_ (.A0(net115),
    .A1(net30),
    .S(net16),
    .X(_0056_));
 sky130_fd_sc_hd__mux2_1 _1042_ (.A0(net117),
    .A1(net28),
    .S(net16),
    .X(_0057_));
 sky130_fd_sc_hd__and4b_2 _1043_ (.A_N(net21),
    .B(_0481_),
    .C(_0485_),
    .D(net22),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_1 _1044_ (.A0(net94),
    .A1(net34),
    .S(_0524_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _1045_ (.A0(net65),
    .A1(net32),
    .S(_0524_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _1046_ (.A0(net98),
    .A1(net30),
    .S(_0524_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _1047_ (.A0(net78),
    .A1(net28),
    .S(_0524_),
    .X(_0061_));
 sky130_fd_sc_hd__and3_2 _1048_ (.A(_0479_),
    .B(_0485_),
    .C(_0514_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_1 _1049_ (.A0(net101),
    .A1(net35),
    .S(_0525_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _1050_ (.A0(net71),
    .A1(net33),
    .S(_0525_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _1051_ (.A0(net106),
    .A1(net31),
    .S(_0525_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _1052_ (.A0(net95),
    .A1(net29),
    .S(_0525_),
    .X(_0065_));
 sky130_fd_sc_hd__nor2_2 _1053_ (.A(_0486_),
    .B(_0516_),
    .Y(_0526_));
 sky130_fd_sc_hd__mux2_1 _1054_ (.A0(net118),
    .A1(net35),
    .S(_0526_),
    .X(_0066_));
 sky130_fd_sc_hd__mux2_1 _1055_ (.A0(net103),
    .A1(net33),
    .S(_0526_),
    .X(_0067_));
 sky130_fd_sc_hd__mux2_1 _1056_ (.A0(net87),
    .A1(net31),
    .S(_0526_),
    .X(_0068_));
 sky130_fd_sc_hd__mux2_1 _1057_ (.A0(net75),
    .A1(net29),
    .S(_0526_),
    .X(_0069_));
 sky130_fd_sc_hd__nor2_2 _1058_ (.A(_0486_),
    .B(_0518_),
    .Y(_0527_));
 sky130_fd_sc_hd__mux2_1 _1059_ (.A0(net79),
    .A1(net35),
    .S(_0527_),
    .X(_0070_));
 sky130_fd_sc_hd__mux2_1 _1060_ (.A0(net77),
    .A1(net33),
    .S(_0527_),
    .X(_0071_));
 sky130_fd_sc_hd__mux2_1 _1061_ (.A0(net73),
    .A1(net31),
    .S(_0527_),
    .X(_0072_));
 sky130_fd_sc_hd__mux2_1 _1062_ (.A0(net99),
    .A1(net29),
    .S(_0527_),
    .X(_0073_));
 sky130_fd_sc_hd__and3_2 _1063_ (.A(_0481_),
    .B(_0485_),
    .C(_0514_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_1 _1064_ (.A0(net84),
    .A1(net35),
    .S(_0528_),
    .X(_0074_));
 sky130_fd_sc_hd__mux2_1 _1065_ (.A0(net104),
    .A1(net33),
    .S(_0528_),
    .X(_0075_));
 sky130_fd_sc_hd__mux2_1 _1066_ (.A0(net85),
    .A1(net31),
    .S(_0528_),
    .X(_0076_));
 sky130_fd_sc_hd__mux2_1 _1067_ (.A0(net74),
    .A1(net29),
    .S(_0528_),
    .X(_0077_));
 sky130_fd_sc_hd__dfrtp_4 _1068_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0005_),
    .RESET_B(net46),
    .Q(\start_seg[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1069_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0006_),
    .RESET_B(net40),
    .Q(\start_seg[1] ));
 sky130_fd_sc_hd__dfrtp_4 _1070_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0007_),
    .RESET_B(net42),
    .Q(\start_seg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1071_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0008_),
    .RESET_B(net45),
    .Q(\start_seg[3] ));
 sky130_fd_sc_hd__dfrtp_4 _1072_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0009_),
    .RESET_B(net46),
    .Q(mode_dec));
 sky130_fd_sc_hd__dfrtp_1 _1073_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0010_),
    .RESET_B(net44),
    .Q(\curr_seg[0] ));
 sky130_fd_sc_hd__dfrtp_1 _1074_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0011_),
    .RESET_B(net44),
    .Q(\curr_seg[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1075_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0012_),
    .RESET_B(net45),
    .Q(\curr_seg[2] ));
 sky130_fd_sc_hd__dfrtp_2 _1076_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0013_),
    .RESET_B(net45),
    .Q(\curr_seg[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1077_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0014_),
    .RESET_B(net43),
    .Q(\full_key[4] ));
 sky130_fd_sc_hd__dfrtp_1 _1078_ (.CLK(clknet_3_6__leaf_clk),
    .D(_0015_),
    .RESET_B(net44),
    .Q(\full_key[5] ));
 sky130_fd_sc_hd__dfrtp_1 _1079_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0016_),
    .RESET_B(net44),
    .Q(\full_key[6] ));
 sky130_fd_sc_hd__dfrtp_1 _1080_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0017_),
    .RESET_B(net43),
    .Q(\full_key[7] ));
 sky130_fd_sc_hd__dfrtp_1 _1081_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0018_),
    .RESET_B(net43),
    .Q(\full_key[12] ));
 sky130_fd_sc_hd__dfrtp_1 _1082_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0019_),
    .RESET_B(net45),
    .Q(\full_key[13] ));
 sky130_fd_sc_hd__dfrtp_1 _1083_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0020_),
    .RESET_B(net44),
    .Q(\full_key[14] ));
 sky130_fd_sc_hd__dfrtp_1 _1084_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0021_),
    .RESET_B(net43),
    .Q(\full_key[15] ));
 sky130_fd_sc_hd__dfrtp_1 _1085_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0022_),
    .RESET_B(net43),
    .Q(\full_key[20] ));
 sky130_fd_sc_hd__dfrtp_1 _1086_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0023_),
    .RESET_B(net44),
    .Q(\full_key[21] ));
 sky130_fd_sc_hd__dfrtp_1 _1087_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0024_),
    .RESET_B(net44),
    .Q(\full_key[22] ));
 sky130_fd_sc_hd__dfrtp_1 _1088_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0025_),
    .RESET_B(net43),
    .Q(\full_key[23] ));
 sky130_fd_sc_hd__dfrtp_1 _1089_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0026_),
    .RESET_B(net43),
    .Q(\full_key[28] ));
 sky130_fd_sc_hd__dfrtp_1 _1090_ (.CLK(clknet_3_7__leaf_clk),
    .D(_0027_),
    .RESET_B(net44),
    .Q(\full_key[29] ));
 sky130_fd_sc_hd__dfrtp_1 _1091_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0028_),
    .RESET_B(net44),
    .Q(\full_key[30] ));
 sky130_fd_sc_hd__dfrtp_1 _1092_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0029_),
    .RESET_B(net43),
    .Q(\full_key[31] ));
 sky130_fd_sc_hd__dfrtp_1 _1093_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0030_),
    .RESET_B(net37),
    .Q(\full_key[36] ));
 sky130_fd_sc_hd__dfrtp_1 _1094_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0031_),
    .RESET_B(net37),
    .Q(\full_key[37] ));
 sky130_fd_sc_hd__dfrtp_1 _1095_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0032_),
    .RESET_B(net37),
    .Q(\full_key[38] ));
 sky130_fd_sc_hd__dfrtp_1 _1096_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0033_),
    .RESET_B(net37),
    .Q(\full_key[39] ));
 sky130_fd_sc_hd__dfrtp_1 _1097_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0034_),
    .RESET_B(net37),
    .Q(\full_key[44] ));
 sky130_fd_sc_hd__dfrtp_1 _1098_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0035_),
    .RESET_B(net37),
    .Q(\full_key[45] ));
 sky130_fd_sc_hd__dfrtp_1 _1099_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0036_),
    .RESET_B(net37),
    .Q(\full_key[46] ));
 sky130_fd_sc_hd__dfrtp_1 _1100_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0037_),
    .RESET_B(net37),
    .Q(\full_key[47] ));
 sky130_fd_sc_hd__dfrtp_1 _1101_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0038_),
    .RESET_B(net37),
    .Q(\full_key[52] ));
 sky130_fd_sc_hd__dfrtp_1 _1102_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0039_),
    .RESET_B(net37),
    .Q(\full_key[53] ));
 sky130_fd_sc_hd__dfrtp_1 _1103_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0040_),
    .RESET_B(net38),
    .Q(\full_key[54] ));
 sky130_fd_sc_hd__dfrtp_1 _1104_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0041_),
    .RESET_B(net38),
    .Q(\full_key[55] ));
 sky130_fd_sc_hd__dfrtp_1 _1105_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0042_),
    .RESET_B(net38),
    .Q(\full_key[60] ));
 sky130_fd_sc_hd__dfrtp_1 _1106_ (.CLK(clknet_3_2__leaf_clk),
    .D(_0043_),
    .RESET_B(net38),
    .Q(\full_key[61] ));
 sky130_fd_sc_hd__dfrtp_1 _1107_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0044_),
    .RESET_B(net40),
    .Q(\full_key[62] ));
 sky130_fd_sc_hd__dfrtp_1 _1108_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0045_),
    .RESET_B(net38),
    .Q(\full_key[63] ));
 sky130_fd_sc_hd__dfrtp_1 _1109_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0046_),
    .RESET_B(net39),
    .Q(\full_key[68] ));
 sky130_fd_sc_hd__dfrtp_1 _1110_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0047_),
    .RESET_B(net39),
    .Q(\full_key[69] ));
 sky130_fd_sc_hd__dfrtp_1 _1111_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0048_),
    .RESET_B(net42),
    .Q(\full_key[70] ));
 sky130_fd_sc_hd__dfrtp_1 _1112_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0049_),
    .RESET_B(net42),
    .Q(\full_key[71] ));
 sky130_fd_sc_hd__dfrtp_1 _1113_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0050_),
    .RESET_B(net39),
    .Q(\full_key[76] ));
 sky130_fd_sc_hd__dfrtp_1 _1114_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0051_),
    .RESET_B(net39),
    .Q(\full_key[77] ));
 sky130_fd_sc_hd__dfrtp_1 _1115_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0052_),
    .RESET_B(net42),
    .Q(\full_key[78] ));
 sky130_fd_sc_hd__dfrtp_1 _1116_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0053_),
    .RESET_B(net42),
    .Q(\full_key[79] ));
 sky130_fd_sc_hd__dfrtp_1 _1117_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0054_),
    .RESET_B(net39),
    .Q(\full_key[84] ));
 sky130_fd_sc_hd__dfrtp_1 _1118_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0055_),
    .RESET_B(net42),
    .Q(\full_key[85] ));
 sky130_fd_sc_hd__dfrtp_1 _1119_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0056_),
    .RESET_B(net42),
    .Q(\full_key[86] ));
 sky130_fd_sc_hd__dfrtp_1 _1120_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0057_),
    .RESET_B(net42),
    .Q(\full_key[87] ));
 sky130_fd_sc_hd__dfrtp_1 _1121_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0058_),
    .RESET_B(net42),
    .Q(\full_key[92] ));
 sky130_fd_sc_hd__dfrtp_1 _1122_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0059_),
    .RESET_B(net42),
    .Q(\full_key[93] ));
 sky130_fd_sc_hd__dfrtp_1 _1123_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0060_),
    .RESET_B(net43),
    .Q(\full_key[94] ));
 sky130_fd_sc_hd__dfrtp_1 _1124_ (.CLK(clknet_3_5__leaf_clk),
    .D(_0061_),
    .RESET_B(net43),
    .Q(\full_key[95] ));
 sky130_fd_sc_hd__dfrtp_1 _1125_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0062_),
    .RESET_B(net39),
    .Q(\full_key[100] ));
 sky130_fd_sc_hd__dfrtp_1 _1126_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0063_),
    .RESET_B(net36),
    .Q(\full_key[101] ));
 sky130_fd_sc_hd__dfrtp_1 _1127_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0064_),
    .RESET_B(net36),
    .Q(\full_key[102] ));
 sky130_fd_sc_hd__dfrtp_1 _1128_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0065_),
    .RESET_B(net36),
    .Q(\full_key[103] ));
 sky130_fd_sc_hd__dfrtp_1 _1129_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0066_),
    .RESET_B(net36),
    .Q(\full_key[108] ));
 sky130_fd_sc_hd__dfrtp_1 _1130_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0067_),
    .RESET_B(net36),
    .Q(\full_key[109] ));
 sky130_fd_sc_hd__dfrtp_1 _1131_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0068_),
    .RESET_B(net36),
    .Q(\full_key[110] ));
 sky130_fd_sc_hd__dfrtp_1 _1132_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0069_),
    .RESET_B(net36),
    .Q(\full_key[111] ));
 sky130_fd_sc_hd__dfrtp_1 _1133_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0070_),
    .RESET_B(net39),
    .Q(\full_key[116] ));
 sky130_fd_sc_hd__dfrtp_1 _1134_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0071_),
    .RESET_B(net36),
    .Q(\full_key[117] ));
 sky130_fd_sc_hd__dfrtp_1 _1135_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0072_),
    .RESET_B(net39),
    .Q(\full_key[118] ));
 sky130_fd_sc_hd__dfrtp_1 _1136_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0073_),
    .RESET_B(net36),
    .Q(\full_key[119] ));
 sky130_fd_sc_hd__dfrtp_1 _1137_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0074_),
    .RESET_B(net39),
    .Q(\full_key[124] ));
 sky130_fd_sc_hd__dfrtp_1 _1138_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0075_),
    .RESET_B(net36),
    .Q(\full_key[125] ));
 sky130_fd_sc_hd__dfrtp_1 _1139_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0076_),
    .RESET_B(net39),
    .Q(\full_key[126] ));
 sky130_fd_sc_hd__dfrtp_1 _1140_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0077_),
    .RESET_B(net41),
    .Q(\full_key[127] ));
 sky130_fd_sc_hd__dfrtp_4 _1141_ (.CLK(clknet_3_3__leaf_clk),
    .D(_0000_),
    .RESET_B(net40),
    .Q(\counter[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1142_ (.CLK(clknet_3_0__leaf_clk),
    .D(_0001_),
    .RESET_B(net38),
    .Q(\counter[1] ));
 sky130_fd_sc_hd__dfrtp_1 _1143_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0002_),
    .RESET_B(net40),
    .Q(\counter[2] ));
 sky130_fd_sc_hd__dfrtp_1 _1144_ (.CLK(clknet_3_1__leaf_clk),
    .D(_0003_),
    .RESET_B(net40),
    .Q(\counter[3] ));
 sky130_fd_sc_hd__dfrtp_1 _1145_ (.CLK(clknet_3_4__leaf_clk),
    .D(_0004_),
    .RESET_B(net40),
    .Q(\counter[4] ));
 sky130_fd_sc_hd__dfrtp_4 _1146_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sys_next_state[0] ),
    .RESET_B(net40),
    .Q(\sys_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _1147_ (.CLK(clknet_3_6__leaf_clk),
    .D(\sys_next_state[1] ),
    .RESET_B(net44),
    .Q(\sys_state[1] ));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_48 (.LO(net48));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_49 (.LO(net49));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_50 (.LO(net50));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_51 (.LO(net51));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_52 (.LO(net52));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_53 (.LO(net53));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_54 (.LO(net54));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_55 (.LO(net55));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_56 (.LO(net56));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_57 (.LO(net57));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_58 (.LO(net58));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_59 (.LO(net59));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_60 (.LO(net60));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_61 (.LO(net61));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_62 (.LO(net62));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_77 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_78 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_79 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_80 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_81 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_82 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_83 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_84 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_85 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_86 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_87 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_88 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_89 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_90 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_91 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_92 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_93 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_94 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_95 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_96 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_97 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_98 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_302 ();
 sky130_fd_sc_hd__clkbuf_1 input1 (.A(rst_n),
    .X(net1));
 sky130_fd_sc_hd__buf_2 input2 (.A(ui_in[0]),
    .X(net2));
 sky130_fd_sc_hd__buf_2 input3 (.A(ui_in[1]),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(ui_in[2]),
    .X(net4));
 sky130_fd_sc_hd__clkbuf_2 input5 (.A(ui_in[3]),
    .X(net5));
 sky130_fd_sc_hd__buf_1 input6 (.A(ui_in[4]),
    .X(net6));
 sky130_fd_sc_hd__dlymetal6s2s_1 input7 (.A(ui_in[5]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(ui_in[6]),
    .X(net8));
 sky130_fd_sc_hd__buf_1 input9 (.A(ui_in[7]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(uio_in[0]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(uio_in[1]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_4 fanout12 (.A(_0143_),
    .X(net12));
 sky130_fd_sc_hd__buf_2 fanout13 (.A(net14),
    .X(net13));
 sky130_fd_sc_hd__buf_2 fanout14 (.A(_0142_),
    .X(net14));
 sky130_fd_sc_hd__buf_2 fanout15 (.A(_0125_),
    .X(net15));
 sky130_fd_sc_hd__buf_1 max_cap16 (.A(net17),
    .X(net16));
 sky130_fd_sc_hd__buf_1 wire17 (.A(_0523_),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_4 fanout18 (.A(net19),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_4 fanout19 (.A(_0085_),
    .X(net19));
 sky130_fd_sc_hd__buf_2 fanout20 (.A(\sys_state[1] ),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 fanout21 (.A(\counter[4] ),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 fanout22 (.A(\counter[2] ),
    .X(net22));
 sky130_fd_sc_hd__buf_2 fanout23 (.A(\curr_seg[2] ),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_4 fanout24 (.A(\curr_seg[1] ),
    .X(net24));
 sky130_fd_sc_hd__buf_2 fanout25 (.A(\curr_seg[1] ),
    .X(net25));
 sky130_fd_sc_hd__buf_4 fanout26 (.A(\curr_seg[0] ),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_4 fanout27 (.A(\curr_seg[0] ),
    .X(net27));
 sky130_fd_sc_hd__clkbuf_4 fanout28 (.A(net29),
    .X(net28));
 sky130_fd_sc_hd__buf_2 fanout29 (.A(net9),
    .X(net29));
 sky130_fd_sc_hd__buf_2 fanout30 (.A(net31),
    .X(net30));
 sky130_fd_sc_hd__buf_2 fanout31 (.A(net8),
    .X(net31));
 sky130_fd_sc_hd__buf_2 fanout32 (.A(net33),
    .X(net32));
 sky130_fd_sc_hd__buf_2 fanout33 (.A(net7),
    .X(net33));
 sky130_fd_sc_hd__buf_2 fanout34 (.A(net35),
    .X(net34));
 sky130_fd_sc_hd__buf_2 fanout35 (.A(net6),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_4 fanout36 (.A(net41),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_4 fanout37 (.A(net41),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 fanout38 (.A(net41),
    .X(net38));
 sky130_fd_sc_hd__clkbuf_4 fanout39 (.A(net41),
    .X(net39));
 sky130_fd_sc_hd__buf_2 fanout40 (.A(net41),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 fanout41 (.A(net46),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_4 fanout42 (.A(net45),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_4 fanout43 (.A(net45),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_4 fanout44 (.A(net45),
    .X(net44));
 sky130_fd_sc_hd__buf_2 fanout45 (.A(net46),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 fanout46 (.A(net1),
    .X(net46));
 sky130_fd_sc_hd__conb_1 tt_um_Samcooper01_47 (.LO(net47));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__bufinv_16 clkload0 (.A(clknet_3_1__leaf_clk));
 sky130_fd_sc_hd__clkinvlp_4 clkload1 (.A(clknet_3_2__leaf_clk));
 sky130_fd_sc_hd__inv_6 clkload2 (.A(clknet_3_3__leaf_clk));
 sky130_fd_sc_hd__clkinv_2 clkload3 (.A(clknet_3_4__leaf_clk));
 sky130_fd_sc_hd__clkbuf_4 clkload4 (.A(clknet_3_5__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload5 (.A(clknet_3_6__leaf_clk));
 sky130_fd_sc_hd__clkinv_4 clkload6 (.A(clknet_3_7__leaf_clk));
 sky130_fd_sc_hd__dlygate4sd3_1 hold1 (.A(\full_key[55] ),
    .X(net63));
 sky130_fd_sc_hd__dlygate4sd3_1 hold2 (.A(\full_key[53] ),
    .X(net64));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(\full_key[93] ),
    .X(net65));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(\full_key[78] ),
    .X(net66));
 sky130_fd_sc_hd__dlygate4sd3_1 hold5 (.A(\full_key[52] ),
    .X(net67));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(\full_key[79] ),
    .X(net68));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(\full_key[54] ),
    .X(net69));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(\full_key[84] ),
    .X(net70));
 sky130_fd_sc_hd__dlygate4sd3_1 hold9 (.A(\full_key[101] ),
    .X(net71));
 sky130_fd_sc_hd__dlygate4sd3_1 hold10 (.A(\full_key[63] ),
    .X(net72));
 sky130_fd_sc_hd__dlygate4sd3_1 hold11 (.A(\full_key[118] ),
    .X(net73));
 sky130_fd_sc_hd__dlygate4sd3_1 hold12 (.A(\full_key[127] ),
    .X(net74));
 sky130_fd_sc_hd__dlygate4sd3_1 hold13 (.A(\full_key[111] ),
    .X(net75));
 sky130_fd_sc_hd__dlygate4sd3_1 hold14 (.A(\full_key[46] ),
    .X(net76));
 sky130_fd_sc_hd__dlygate4sd3_1 hold15 (.A(\full_key[117] ),
    .X(net77));
 sky130_fd_sc_hd__dlygate4sd3_1 hold16 (.A(\full_key[95] ),
    .X(net78));
 sky130_fd_sc_hd__dlygate4sd3_1 hold17 (.A(\full_key[116] ),
    .X(net79));
 sky130_fd_sc_hd__dlygate4sd3_1 hold18 (.A(\full_key[60] ),
    .X(net80));
 sky130_fd_sc_hd__dlygate4sd3_1 hold19 (.A(\full_key[62] ),
    .X(net81));
 sky130_fd_sc_hd__dlygate4sd3_1 hold20 (.A(\full_key[29] ),
    .X(net82));
 sky130_fd_sc_hd__dlygate4sd3_1 hold21 (.A(\full_key[30] ),
    .X(net83));
 sky130_fd_sc_hd__dlygate4sd3_1 hold22 (.A(\full_key[124] ),
    .X(net84));
 sky130_fd_sc_hd__dlygate4sd3_1 hold23 (.A(\full_key[126] ),
    .X(net85));
 sky130_fd_sc_hd__dlygate4sd3_1 hold24 (.A(\full_key[61] ),
    .X(net86));
 sky130_fd_sc_hd__dlygate4sd3_1 hold25 (.A(\full_key[110] ),
    .X(net87));
 sky130_fd_sc_hd__dlygate4sd3_1 hold26 (.A(\full_key[28] ),
    .X(net88));
 sky130_fd_sc_hd__dlygate4sd3_1 hold27 (.A(\full_key[6] ),
    .X(net89));
 sky130_fd_sc_hd__dlygate4sd3_1 hold28 (.A(\full_key[15] ),
    .X(net90));
 sky130_fd_sc_hd__dlygate4sd3_1 hold29 (.A(\full_key[22] ),
    .X(net91));
 sky130_fd_sc_hd__dlygate4sd3_1 hold30 (.A(\full_key[5] ),
    .X(net92));
 sky130_fd_sc_hd__dlygate4sd3_1 hold31 (.A(\full_key[85] ),
    .X(net93));
 sky130_fd_sc_hd__dlygate4sd3_1 hold32 (.A(\full_key[92] ),
    .X(net94));
 sky130_fd_sc_hd__dlygate4sd3_1 hold33 (.A(\full_key[103] ),
    .X(net95));
 sky130_fd_sc_hd__dlygate4sd3_1 hold34 (.A(\full_key[71] ),
    .X(net96));
 sky130_fd_sc_hd__dlygate4sd3_1 hold35 (.A(\full_key[70] ),
    .X(net97));
 sky130_fd_sc_hd__dlygate4sd3_1 hold36 (.A(\full_key[94] ),
    .X(net98));
 sky130_fd_sc_hd__dlygate4sd3_1 hold37 (.A(\full_key[119] ),
    .X(net99));
 sky130_fd_sc_hd__dlygate4sd3_1 hold38 (.A(\full_key[14] ),
    .X(net100));
 sky130_fd_sc_hd__dlygate4sd3_1 hold39 (.A(\full_key[100] ),
    .X(net101));
 sky130_fd_sc_hd__dlygate4sd3_1 hold40 (.A(\full_key[4] ),
    .X(net102));
 sky130_fd_sc_hd__dlygate4sd3_1 hold41 (.A(\full_key[109] ),
    .X(net103));
 sky130_fd_sc_hd__dlygate4sd3_1 hold42 (.A(\full_key[125] ),
    .X(net104));
 sky130_fd_sc_hd__dlygate4sd3_1 hold43 (.A(\full_key[23] ),
    .X(net105));
 sky130_fd_sc_hd__dlygate4sd3_1 hold44 (.A(\full_key[102] ),
    .X(net106));
 sky130_fd_sc_hd__dlygate4sd3_1 hold45 (.A(\full_key[76] ),
    .X(net107));
 sky130_fd_sc_hd__dlygate4sd3_1 hold46 (.A(\full_key[69] ),
    .X(net108));
 sky130_fd_sc_hd__dlygate4sd3_1 hold47 (.A(\full_key[37] ),
    .X(net109));
 sky130_fd_sc_hd__dlygate4sd3_1 hold48 (.A(\full_key[31] ),
    .X(net110));
 sky130_fd_sc_hd__dlygate4sd3_1 hold49 (.A(\full_key[45] ),
    .X(net111));
 sky130_fd_sc_hd__dlygate4sd3_1 hold50 (.A(\full_key[77] ),
    .X(net112));
 sky130_fd_sc_hd__dlygate4sd3_1 hold51 (.A(\full_key[68] ),
    .X(net113));
 sky130_fd_sc_hd__dlygate4sd3_1 hold52 (.A(\full_key[12] ),
    .X(net114));
 sky130_fd_sc_hd__dlygate4sd3_1 hold53 (.A(\full_key[86] ),
    .X(net115));
 sky130_fd_sc_hd__dlygate4sd3_1 hold54 (.A(\full_key[47] ),
    .X(net116));
 sky130_fd_sc_hd__dlygate4sd3_1 hold55 (.A(\full_key[87] ),
    .X(net117));
 sky130_fd_sc_hd__dlygate4sd3_1 hold56 (.A(\full_key[108] ),
    .X(net118));
 sky130_fd_sc_hd__dlygate4sd3_1 hold57 (.A(\full_key[39] ),
    .X(net119));
 sky130_fd_sc_hd__dlygate4sd3_1 hold58 (.A(\full_key[21] ),
    .X(net120));
 sky130_fd_sc_hd__dlygate4sd3_1 hold59 (.A(\full_key[13] ),
    .X(net121));
 sky130_fd_sc_hd__dlygate4sd3_1 hold60 (.A(\full_key[7] ),
    .X(net122));
 sky130_fd_sc_hd__dlygate4sd3_1 hold61 (.A(\full_key[20] ),
    .X(net123));
 sky130_fd_sc_hd__dlygate4sd3_1 hold62 (.A(\full_key[36] ),
    .X(net124));
 sky130_fd_sc_hd__dlygate4sd3_1 hold63 (.A(\full_key[38] ),
    .X(net125));
 sky130_fd_sc_hd__dlygate4sd3_1 hold64 (.A(\full_key[44] ),
    .X(net126));
 sky130_fd_sc_hd__dlygate4sd3_1 hold65 (.A(\counter[0] ),
    .X(net127));
 sky130_ef_sc_hd__decap_12 FILLER_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_192 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_87 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_1_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_1_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_1_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_1_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_1_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_1_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_137 ();
 sky130_fd_sc_hd__decap_4 FILLER_2_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_2_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_2_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_2_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_2_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_2_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_2_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_106 ();
 sky130_fd_sc_hd__decap_3 FILLER_3_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_3_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_3_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_3_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_3_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_3_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_91 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_4_217 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_4_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_4_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_290 ();
 sky130_fd_sc_hd__decap_6 FILLER_4_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_4_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_4_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_122 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_147 ();
 sky130_fd_sc_hd__decap_8 FILLER_5_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_5_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_212 ();
 sky130_fd_sc_hd__decap_6 FILLER_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_5_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_5_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_5_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_119 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_150 ();
 sky130_fd_sc_hd__decap_3 FILLER_6_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_6_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_6_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_259 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_6_297 ();
 sky130_fd_sc_hd__decap_8 FILLER_6_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_6_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_223 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_7_252 ();
 sky130_fd_sc_hd__fill_2 FILLER_7_278 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_7_294 ();
 sky130_fd_sc_hd__decap_4 FILLER_7_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_7_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_8_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_94 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_8_214 ();
 sky130_fd_sc_hd__decap_3 FILLER_8_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_8_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_8_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_8_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_9_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_9_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_9_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_9_252 ();
 sky130_fd_sc_hd__decap_4 FILLER_9_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_9_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_296 ();
 sky130_fd_sc_hd__fill_1 FILLER_9_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_10_212 ();
 sky130_fd_sc_hd__decap_8 FILLER_10_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_238 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_10_257 ();
 sky130_fd_sc_hd__fill_2 FILLER_10_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_10_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_11_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_35 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_11_104 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_11_201 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_11_274 ();
 sky130_fd_sc_hd__decap_3 FILLER_11_289 ();
 sky130_fd_sc_hd__fill_2 FILLER_11_301 ();
 sky130_fd_sc_hd__decap_4 FILLER_11_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_158 ();
 sky130_fd_sc_hd__decap_3 FILLER_12_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_12_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_12_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_12_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_12_282 ();
 sky130_fd_sc_hd__decap_4 FILLER_12_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_12_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_13_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_179 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_13_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_13_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_13_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_13_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_13_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_146 ();
 sky130_fd_sc_hd__decap_3 FILLER_14_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_14_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_14_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_14_326 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_147 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_173 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_15_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_236 ();
 sky130_fd_sc_hd__decap_8 FILLER_15_248 ();
 sky130_fd_sc_hd__decap_3 FILLER_15_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_15_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_285 ();
 sky130_fd_sc_hd__decap_4 FILLER_15_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_15_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_15_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_16_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_108 ();
 sky130_fd_sc_hd__decap_8 FILLER_16_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_16_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_16_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_16_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_16_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_16_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_17_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_212 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_17_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_17_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_17_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_17_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_49 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_98 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_18_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_18_195 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_261 ();
 sky130_fd_sc_hd__decap_3 FILLER_18_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_18_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_18_325 ();
 sky130_fd_sc_hd__fill_2 FILLER_18_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_19_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_208 ();
 sky130_fd_sc_hd__decap_8 FILLER_19_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_19_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_19_239 ();
 sky130_fd_sc_hd__fill_2 FILLER_19_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_19_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_19_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_105 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_117 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_153 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_165 ();
 sky130_fd_sc_hd__decap_3 FILLER_20_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_246 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_266 ();
 sky130_fd_sc_hd__decap_6 FILLER_20_278 ();
 sky130_fd_sc_hd__fill_1 FILLER_20_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_20_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_20_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_21_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_21_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_21_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_21_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_21_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_92 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_22_176 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_226 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_22_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_250 ();
 sky130_fd_sc_hd__fill_2 FILLER_22_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_280 ();
 sky130_fd_sc_hd__decap_6 FILLER_22_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_22_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_22_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_22_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_98 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_130 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_142 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_174 ();
 sky130_fd_sc_hd__decap_6 FILLER_23_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_23_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_235 ();
 sky130_fd_sc_hd__decap_8 FILLER_23_247 ();
 sky130_fd_sc_hd__decap_3 FILLER_23_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_23_293 ();
 sky130_fd_sc_hd__decap_4 FILLER_23_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_118 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_24_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_24_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_227 ();
 sky130_fd_sc_hd__fill_2 FILLER_24_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_240 ();
 sky130_ef_sc_hd__decap_12 FILLER_24_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_24_292 ();
 sky130_fd_sc_hd__decap_3 FILLER_24_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_24_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_87 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_95 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_25_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_248 ();
 sky130_fd_sc_hd__decap_6 FILLER_25_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_25_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_25_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_25_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_25_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_25_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_45 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_26_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_200 ();
 sky130_fd_sc_hd__decap_8 FILLER_26_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_26_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_26_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_26_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_26_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_26_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_94 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_118 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_27_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_257 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_27_288 ();
 sky130_fd_sc_hd__fill_2 FILLER_27_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_27_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_27_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_27_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_48 ();
 sky130_fd_sc_hd__decap_6 FILLER_28_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_66 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_132 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_159 ();
 sky130_fd_sc_hd__decap_4 FILLER_28_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_280 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_292 ();
 sky130_fd_sc_hd__fill_2 FILLER_28_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_28_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_28_312 ();
 sky130_fd_sc_hd__decap_8 FILLER_28_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_28_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_200 ();
 sky130_fd_sc_hd__decap_3 FILLER_29_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_229 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_234 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_29_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_29_289 ();
 sky130_fd_sc_hd__fill_1 FILLER_29_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_29_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_29_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_56 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_112 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_152 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_30_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_30_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_30_287 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_30_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_30_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_31_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_31_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_31_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_31_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_31_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_31_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_104 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_116 ();
 sky130_fd_sc_hd__fill_2 FILLER_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_32_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_205 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_32_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_32_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_32_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_32_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_33_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_235 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_33_267 ();
 sky130_fd_sc_hd__decap_4 FILLER_33_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_33_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_33_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_33_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_34_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_211 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_34_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_34_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_34_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_34_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_34_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_34_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_147 ();
 sky130_fd_sc_hd__decap_4 FILLER_35_159 ();
 sky130_fd_sc_hd__fill_2 FILLER_35_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_35_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_35_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_35_299 ();
 sky130_fd_sc_hd__decap_3 FILLER_35_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_35_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_144 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_36_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_36_302 ();
 sky130_fd_sc_hd__decap_4 FILLER_36_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_36_326 ();
 sky130_fd_sc_hd__fill_1 FILLER_36_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_37_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_37_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_155 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_37_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_37_248 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_291 ();
 sky130_fd_sc_hd__decap_3 FILLER_37_303 ();
 sky130_ef_sc_hd__decap_12 FILLER_37_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_37_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_70 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_88 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_94 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_100 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_124 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_130 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_136 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_148 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_160 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_38_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_38_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_38_299 ();
 sky130_fd_sc_hd__decap_4 FILLER_38_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_38_316 ();
 sky130_fd_sc_hd__decap_6 FILLER_38_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_38_334 ();
 assign uio_oe[0] = net47;
 assign uio_oe[1] = net48;
 assign uio_oe[2] = net49;
 assign uio_oe[3] = net50;
 assign uio_oe[4] = net51;
 assign uio_oe[5] = net52;
 assign uio_oe[6] = net53;
 assign uio_oe[7] = net54;
 assign uio_out[0] = net55;
 assign uio_out[1] = net56;
 assign uio_out[2] = net57;
 assign uio_out[3] = net58;
 assign uio_out[4] = net59;
 assign uio_out[5] = net60;
 assign uio_out[6] = net61;
 assign uio_out[7] = net62;
endmodule
